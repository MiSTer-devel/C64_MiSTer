
module sid_filters
#(
	parameter MULTI_FILTERS = 1
)
(
	input             clk,
	input             rst,
	input      [10:0] Fc,
	input       [7:0] Res_Filt,
	input       [7:0] Mode_Vol,
	input      [17:0] voice1,
	input      [17:0] voice2,
	input      [17:0] voice3,
	input      [17:0] ext_in,
	input             input_valid,
	input             enable,
	output reg [17:0] sound,

	input             mode,
	input       [1:0] mixctl,
	input       [2:0] cfg,
	input             ld_clk,
	input      [11:0] ld_addr,
	input      [15:0] ld_data,
	input             ld_wr
);

reg signed [17:0] Vhp;
reg signed [17:0] Vbp;
reg signed [17:0] w0;
reg signed [17:0] q;

wire [10:0] divmul[32] =
'{
	1448, 1323, 1218, 1128, 1051, 984, 925, 872,
	 825,  783,  745,  710,  679, 650, 624, 599,
	 
	1448, 1328, 1218, 1117, 1024, 939, 861, 790,
	 724,  664,  609,  558,  512, 470, 431, 395
};

wire [35:0] mul1 = w0 * Vhp;
wire [35:0] mul2 = w0 * Vbp;
wire [35:0] mul3 = q  * Vbp;
wire [35:0] mul4 = 18'd82355 * (Fc + 1'b1);

function [17:0] add_limit;
	input [17:0] a,b;
begin
	reg [18:0] tmp;
	tmp = {a[17],a} + {b[17],b};
	add_limit = ^tmp[18:17] ? {tmp[18], {17{tmp[17]}}} : tmp[17:0];
end
endfunction

function [17:0] sub_limit;
	input [17:0] a,b;
begin
	reg [18:0] tmp;
	tmp = {a[17],a} - {b[17],b};
	sub_limit = ^tmp[18:17] ? {tmp[18], {17{tmp[17]}}} : tmp[17:0];
end
endfunction

// Filter
always @(posedge clk) begin
	reg [17:0] dVbp;
	reg [17:0] Vlp;
	reg [17:0] dVlp;
	reg [17:0] Vi;
	reg [17:0] Vnf;
	reg [17:0] Vf;
	reg  [3:0] state;
	reg signed [35:0] mulr;
	reg signed [17:0] mula;
	reg signed [17:0] mulb;

	if (rst) begin
		state <= 0;
		Vlp   <= 0;
		Vbp   <= 0;
		Vhp   <= 0;
	end
	else begin
		state <= state + 1'd1;
		case (state)
			0:	if (input_valid) begin
					sound <= ^mulr[21:20] ? {mulr[21], {17{mulr[20]}}} : mulr[20:3];
					Vi    <= 0;
					Vnf   <= 16384;
					Vf    <= 0;
					w0    <= mode ? {mul4[35], mul4[28:12]} : {1'b0, f0, 1'b0};
				end
				else begin
					state <= 0;
				end
			1:	begin
					if(Res_Filt[0])       Vi   <= add_limit(Vi,  voice1);
					else                  Vnf  <= add_limit(Vnf, voice1);
				end
			2:	begin
					if(Res_Filt[1])       Vi   <= add_limit(Vi,  voice2);
					else                  Vnf  <= add_limit(Vnf, voice2);
				end
			3:	begin
					if(Res_Filt[2])       Vi   <= add_limit(Vi,  voice3);
					else if(!Mode_Vol[7]) Vnf  <= add_limit(Vnf, voice3);

					                      dVbp <= {mul1[35], mul1[35:19]}; // w0 * Vhp
				end
			4:	begin
					if(Res_Filt[3])       Vi   <= add_limit(Vi,  ext_in);
					else                  Vnf  <= add_limit(Vnf, ext_in);

					                      dVlp <= {mul2[35], mul2[35:19]}; // w0 * Vbp
					                      Vbp  <= sub_limit(Vbp, dVbp);
					                      q    <= divmul[{mode, Res_Filt[7:4]}];
				end
			5:	begin
					if(Mode_Vol[5])       Vf   <= add_limit(Vf, Vbp);

					                      Vlp  <= sub_limit(Vlp, dVlp);
				end
			6: begin
					if(Mode_Vol[4])       Vf   <= add_limit(Vf, Vlp);

					                      Vhp  <= sub_limit({mul3[35], mul3[26:10]}, Vlp); // q * Vbp
				end
			7: begin
					                      Vhp  <= sub_limit(Vhp, Vi);
				end
			8:	begin
					if(Mode_Vol[6])       Vf   <= add_limit(Vf, Vhp);
				end
			9:	begin
					mula  <= add_limit((mixctl[1] ? 18'd0 : Vnf), enable ? (mixctl[0] ? 18'd0 : mode ? Vf : (Vf - {Vf[17],Vf[17],Vf[17:2]})) : Vi);
					mulb  <= Mode_Vol[3:0];
				end
			10:begin
					mulr  <= mula * mulb;
					state <= 0;
				end
		endcase
	end
end

reg [15:0] f0;
generate
	if(MULTI_FILTERS) begin
		always @(posedge ld_clk) if(ld_wr) f6581_curve[1024+ld_addr] <= ld_data;
		always @(posedge clk) f0 <= f6581_curve[{cfg, Fc[10:1]}];
	end
	else begin
		always @(posedge ld_clk) if(ld_wr) f6581_curve[ld_addr[9:0]] <= ld_data;
		always @(posedge clk) f0 <= f6581_curve[Fc[10:1]];
	end
endgenerate

// value = pi * 1.048576 * f0[fc]
reg  [15:0] f6581_curve[4*1024] =
'{
	// 0 mixed calc 
      933,    932,    932,    933,    936,    937,    943,    948,
      949,    945,    936,    926,    920,    918,    920,    924,
      930,    938,    945,    954,    960,    960,    955,    951,
      950,    949,    948,    948,    948,    945,    945,    945,
      948,    943,    942,    937,    937,    937,    939,    945,
      950,    951,    956,    960,    965,    971,    977,    981,
      982,    979,    976,    970,    964,    957,    949,    944,
      942,    942,    945,    950,    955,    955,    957,    960,
      961,    957,    954,    948,    948,    949,    955,    958,
      964,    971,    975,    979,    981,    979,    979,    975,
      973,    971,    970,    969,    969,    969,    969,    973,
      973,    971,    967,    965,    965,    963,    963,    967,
      970,    976,    987,    995,   1001,    996,    993,    987,
      983,    982,    984,    988,    992,    992,    994,    999,
      999,    994,    988,    981,    982,    988,   1002,   1014,
     1020,   1018,   1008,   1000,    994,    996,    997,   1005,
     1009,   1008,   1006,   1002,   1005,   1006,   1012,   1018,
     1024,   1024,   1024,   1024,   1026,   1027,   1029,   1033,
     1035,   1033,   1029,   1026,   1027,   1029,   1035,   1041,
     1047,   1048,   1047,   1048,   1053,   1059,   1072,   1082,
     1086,   1078,   1063,   1047,   1041,   1045,   1057,   1069,
     1078,   1082,   1086,   1087,   1090,   1090,   1089,   1087,
     1090,   1091,   1098,   1104,   1105,   1099,   1092,   1086,
     1086,   1096,   1115,   1132,   1147,   1150,   1147,   1141,
     1141,   1141,   1144,   1149,   1154,   1156,   1162,   1166,
     1174,   1180,   1187,   1194,   1197,   1193,   1189,   1183,
     1183,   1188,   1197,   1209,   1216,   1216,   1213,   1210,
     1210,   1210,   1213,   1216,   1219,   1220,   1222,   1225,
     1231,   1238,   1247,   1259,   1271,   1275,   1280,   1286,
     1293,   1297,   1303,   1306,   1310,   1308,   1306,   1306,
     1310,   1318,   1330,   1343,   1354,   1360,   1364,   1367,
     1378,   1393,   1415,   1435,   1448,   1448,   1436,   1426,
     1426,   1435,   1451,   1471,   1484,   1486,   1486,   1486,
     1490,   1498,   1510,   1520,   1535,   1545,   1555,   1564,
     1576,   1585,   1599,   1612,   1622,   1625,   1630,   1633,
     1644,   1655,   1676,   1696,   1713,   1723,   1732,   1738,
     1750,   1761,   1777,   1794,   1807,   1818,   1823,   1828,
     1840,   1857,   1880,   1904,   1921,   1931,   1937,   1944,
     1956,   1970,   1992,   2013,   2035,   2053,   2069,   2087,
     2106,   2124,   2145,   2164,   2185,   2204,   2220,   2238,
     2262,   2283,   2308,   2333,   2356,   2375,   2392,   2409,
     2429,   2448,   2468,   2488,   2510,   2537,   2567,   2601,
     2629,   2650,   2672,   2693,   2720,   2757,   2799,   2843,
     2881,   2905,   2927,   2943,   2969,   2993,   3023,   3054,
     3086,   3115,   3145,   3175,   3207,   3243,   3280,   3319,
     3353,   3385,   3415,   3444,   3472,   3493,   3511,   3531,
     3563,   3606,   3660,   3715,   3761,   3787,   3804,   3819,
     3845,   3888,   3941,   3991,   4033,   4051,   4062,   4071,
     4092,   4126,   4169,   4218,   4264,   4303,   4345,   4383,
     4424,   4460,   4493,   4530,   4575,   4629,   4692,   4755,
     4814,   4862,   4903,   4945,   4991,   5045,   5102,   5160,
     5217,   5269,   5316,   5366,   5421,   5480,   5542,   5604,
     5664,   5716,   5763,   5813,   5867,   5929,   5996,   6064,
     6129,   6185,   6240,   6294,   6354,   6415,   6483,   6548,
     6614,   6670,   6723,   6778,   6840,   6910,   6988,   7067,
     7144,   7216,   7287,   7354,   7420,   7481,   7536,   7593,
     7654,   7715,   7777,   7845,   7917,   7996,   8083,   8171,
     8255,   8332,   8408,   8482,   8558,   8628,   8696,   8768,
     8851,   8946,   9057,   9164,   9261,   9336,   9400,   9466,
     9541,   9629,   9727,   9825,   9922,  10011,  10096,  10181,
    10275,  10377,  10485,  10595,  10701,  10789,  10868,  10952,
    11056,  11187,  11336,  11485,  11617,  11719,  11803,  11886,
    11983,  12099,  12228,  12360,  12487,  12601,  12712,  12829,
    12961,  13151,  13389,  13597,  13706,  13649,  13479,  13308,
    10866,  10883,  10985,  11125,  11250,  11362,  11483,  11606,
    11720,  11813,  11899,  11984,  12076,  12180,  12294,  12408,
    12516,  12607,  12689,  12773,  12869,  12976,  13091,  13212,
    13332,  13454,  13578,  13699,  13812,  13911,  14003,  14089,
    14180,  14270,  14362,  14456,  14559,  14666,  14787,  14904,
    15011,  15096,  15172,  15250,  15344,  15458,  15590,  15723,
    15851,  15960,  16063,  16168,  16281,  16408,  16544,  16680,
    16801,  16904,  16995,  17080,  17157,  17216,  17264,  17317,
    17396,  17508,  17647,  17789,  17919,  18027,  18124,  18219,
    18315,  18410,  18504,  18601,  18705,  18821,  18944,  19070,
    19194,  19312,  19431,  19546,  19659,  19762,  19859,  19959,
    20066,  20187,  20318,  20447,  20568,  20669,  20764,  20856,
    20952,  21048,  21147,  21249,  21357,  21470,  21588,  21707,
    21828,  21951,  22076,  22197,  22316,  22424,  22528,  22631,
    22743,  22864,  22992,  23120,  23247,  23367,  23484,  23602,
    23725,  23869,  24031,  24170,  24251,  24230,  24142,  24052,
    24037,  24125,  24274,  24443,  24594,  24714,  24827,  24937,
    25049,  25168,  25289,  25406,  25517,  25609,  25693,  25777,
    25879,  26004,  26147,  26290,  26416,  26514,  26599,  26682,
    26781,  26908,  27050,  27190,  27308,  27392,  27454,  27517,
    27599,  27712,  27845,  27978,  28094,  28181,  28248,  28319,
    28412,  28541,  28691,  28841,  28968,  29059,  29133,  29201,
    29281,  29375,  29476,  29582,  29688,  29797,  29910,  30022,
    30130,  30229,  30326,  30419,  30505,  30578,  30643,  30707,
    30781,  30867,  30960,  31056,  31146,  31228,  31308,  31386,
    31467,  31551,  31635,  31722,  31813,  31904,  31998,  32093,
    32192,  32292,  32395,  32496,  32591,  32674,  32750,  32825,
    32911,  33009,  33116,  33222,  33313,  33383,  33440,  33497,
    33566,  33654,  33752,  33851,  33941,  34014,  34078,  34139,
    34205,  34273,  34344,  34415,  34487,  34559,  34632,  34705,
    34773,  34832,  34888,  34942,  35004,  35073,  35146,  35220,
    35292,  35371,  35458,  35526,  35552,  35506,  35408,  35310,
    35265,  35298,  35375,  35468,  35544,  35594,  35636,  35677,
    35727,  35788,  35855,  35922,  35982,  36033,  36079,  36121,
    36159,  36187,  36207,  36231,  36269,  36327,  36399,  36473,
    36540,  36601,  36659,  36710,  36751,  36771,  36778,  36785,
    36806,  36846,  36899,  36954,  37004,  37047,  37088,  37125,
    37157,  37182,  37200,  37218,  37243,  37276,  37312,  37352,
    37390,  37427,  37466,  37504,  37540,  37574,  37607,  37640,
    37672,  37708,  37745,  37780,  37809,  37829,  37843,  37857,
    37874,  37893,  37914,  37937,  37962,  37992,  38024,  38057,
    38090,  38120,  38151,  38181,  38210,  38238,  38267,  38294,
    38318,  38340,  38359,  38378,  38398,  38418,  38438,  38459,
    38480,  38502,  38525,  38548,  38569,  38590,  38609,  38627,
    38646,  38665,  38685,  38704,  38723,  38742,  38761,  38780,
    38798,  38817,  38837,  38855,  38870,  38880,  38887,  38895,
    38905,  38920,  38937,  38954,  38973,  38992,  39013,  39032,
    39047,  39058,  39065,  39070,  39072,  39071,  39066,  39061,
    39061,  39064,  39070,  39079,  39088,  39099,  39112,  39125,
    39136,  39142,  39143,  39145,  39146,  39148,  39149,  39151,
    39152,  39154,  39155,  39156,  39158,  39159,  39160,  39161,
    39163,  39164,  39165,  39166,  39168,  39169,  39170,  39171,
    39172,  39173,  39174,  39175,  39176,  39177,  39178,  39179,
    39180,  39181,  39182,  39183,  39184,  39185,  39186,  39187,
    39188,  39189,  39189,  39190,  39191,  39192,  39193,  39194,
    39194,  39195,  39196,  39197,  39198,  39198,  39199,  39200,
    39201,  39202,  39202,  39203,  39204,  39204,  39205,  39206,
    39207,  39207,  39208,  39209,  39209,  39210,  39210,  39211,
    39212,  39212,  39213,  39213,  39214,  39214,  39215,  39215,
    39216,  39216,  39217,  39217,  39218,  39218,  39219,  39219,
    39220,  39220,  39220,  39221,  39221,  39222,  39222,  39222,
    39223,  39223,  39224,  39224,  39224,  39225,  39225,  39226,
    39226,  39226,  39227,  39227,  39227,  39228,  39228,  39228,
    39229,  39229,  39229,  39230,  39230,  39231,  39231,  39231,
	 

	// 1 web 
      843,    840,    840,    843,    846,    849,    859,    866,
      869,    859,    843,    826,    816,    813,    816,    823,
      833,    843,    856,    869,    879,    879,    872,    866,
      863,    859,    856,    856,    856,    853,    853,    853,
      853,    846,    843,    836,    836,    836,    840,    846,
      853,    856,    863,    869,    879,    886,    896,    902,
      905,    899,    892,    882,    872,    859,    846,    833,
      830,    830,    836,    843,    849,    849,    853,    856,
      856,    849,    843,    833,    833,    833,    843,    849,
      859,    866,    872,    879,    882,    879,    876,    869,
      866,    863,    859,    856,    856,    856,    856,    859,
      859,    856,    849,    843,    843,    840,    840,    843,
      849,    859,    872,    886,    896,    889,    879,    869,
      863,    859,    863,    869,    872,    872,    876,    879,
      879,    869,    859,    846,    846,    856,    876,    896,
      905,    899,    882,    866,    856,    856,    859,    866,
      872,    869,    863,    856,    856,    859,    866,    876,
      882,    882,    879,    879,    879,    879,    882,    886,
      889,    882,    876,    866,    866,    869,    876,    886,
      892,    892,    889,    889,    892,    902,    922,    935,
      942,    925,    896,    869,    856,    859,    876,    896,
      909,    912,    915,    915,    915,    912,    909,    905,
      905,    905,    912,    919,    919,    905,    889,    872,
      869,    882,    912,    938,    958,    958,    948,    935,
      928,    925,    928,    932,    935,    935,    942,    945,
      952,    958,    968,    975,    978,    968,    955,    942,
      938,    942,    955,    968,    978,    975,    965,    955,
      952,    948,    948,    948,    948,    945,    945,    942,
      948,    955,    968,    981,    994,    998,   1001,   1004,
     1008,   1008,   1011,   1011,   1011,   1001,    991,    981,
      981,    988,    998,   1014,   1024,   1024,   1021,   1017,
     1024,   1040,   1067,   1090,   1103,   1090,   1060,   1031,
     1017,   1021,   1037,   1057,   1067,   1060,   1047,   1034,
     1027,   1027,   1034,   1040,   1050,   1054,   1057,   1060,
     1067,   1070,   1080,   1087,   1090,   1083,   1073,   1067,
     1067,   1073,   1093,   1110,   1123,   1123,   1123,   1116,
     1120,   1123,   1133,   1143,   1149,   1146,   1136,   1129,
     1129,   1139,   1156,   1176,   1185,   1182,   1169,   1159,
     1156,   1159,   1172,   1185,   1199,   1202,   1208,   1212,
     1218,   1222,   1232,   1238,   1245,   1248,   1248,   1251,
     1258,   1264,   1278,   1288,   1297,   1297,   1294,   1291,
     1291,   1288,   1288,   1288,   1294,   1304,   1320,   1340,
     1353,   1353,   1350,   1350,   1360,   1383,   1419,   1456,
     1482,   1485,   1479,   1469,   1469,   1472,   1482,   1492,
     1505,   1512,   1521,   1531,   1544,   1561,   1581,   1604,
     1620,   1630,   1637,   1640,   1643,   1633,   1617,   1604,
     1610,   1640,   1686,   1736,   1765,   1762,   1742,   1719,
     1716,   1739,   1782,   1821,   1841,   1824,   1792,   1755,
     1739,   1745,   1768,   1798,   1821,   1831,   1841,   1848,
     1854,   1851,   1844,   1841,   1851,   1877,   1917,   1956,
     1986,   1996,   1992,   1992,   1999,   2016,   2039,   2062,
     2085,   2095,   2101,   2108,   2124,   2147,   2177,   2207,
     2233,   2243,   2246,   2253,   2266,   2292,   2328,   2365,
     2394,   2411,   2421,   2431,   2447,   2470,   2500,   2529,
     2556,   2566,   2569,   2576,   2595,   2628,   2674,   2724,
     2767,   2800,   2833,   2859,   2882,   2892,   2895,   2898,
     2908,   2918,   2931,   2951,   2981,   3024,   3076,   3136,
     3185,   3221,   3254,   3287,   3317,   3340,   3356,   3379,
     3422,   3491,   3584,   3673,   3742,   3771,   3778,   3785,
     3811,   3860,   3929,   3999,   4065,   4114,   4157,   4200,
     4256,   4328,   4410,   4493,   4562,   4595,   4608,   4628,
     4684,   4793,   4938,   5082,   5194,   5244,   5260,   5270,
     5313,   5395,   5501,   5610,   5708,   5774,   5827,   5886,
     5969,   6143,   6384,   6548,   6506,   6117,   5488,   4849,
     4420,   4282,   4312,   4420,   4516,   4595,   4697,   4802,
     4891,   4941,   4977,   5010,   5059,   5135,   5227,   5320,
     5395,   5438,   5461,   5488,   5534,   5606,   5692,   5791,
     5890,   5992,   6100,   6206,   6295,   6357,   6407,   6450,
     6502,   6558,   6621,   6690,   6776,   6881,   7010,   7135,
     7240,   7303,   7342,   7388,   7467,   7593,   7754,   7919,
     8067,   8182,   8281,   8383,   8505,   8657,   8831,   9003,
     9144,   9246,   9325,   9388,   9437,   9447,   9431,   9427,
     9480,   9615,   9806,  10007,  10182,  10307,  10409,  10505,
    10607,  10706,  10804,  10907,  11032,  11180,  11348,  11523,
    11694,  11852,  12013,  12168,  12317,  12442,  12557,  12676,
    12814,  12985,  13183,  13377,  13549,  13680,  13792,  13898,
    14013,  14135,  14260,  14392,  14540,  14702,  14876,  15057,
    15242,  15430,  15624,  15815,  15996,  16154,  16299,  16444,
    16612,  16803,  17014,  17228,  17439,  17630,  17818,  18006,
    18210,  18473,  18783,  19033,  19129,  18951,  18589,  18226,
    18062,  18174,  18450,  18786,  19070,  19271,  19455,  19633,
    19817,  20018,  20229,  20433,  20615,  20750,  20858,  20970,
    21132,  21362,  21646,  21929,  22166,  22324,  22443,  22558,
    22723,  22967,  23260,  23550,  23777,  23899,  23958,  24018,
    24139,  24357,  24634,  24917,  25147,  25286,  25368,  25460,
    25625,  25902,  26251,  26603,  26883,  27051,  27160,  27256,
    27387,  27569,  27773,  27997,  28224,  28461,  28715,  28969,
    29206,  29423,  29631,  29825,  29996,  30125,  30227,  30326,
    30461,  30639,  30846,  31064,  31261,  31429,  31588,  31746,
    31914,  32092,  32276,  32470,  32678,  32892,  33119,  33353,
    33597,  33854,  34124,  34391,  34635,  34832,  35004,  35178,
    35389,  35659,  35972,  36279,  36532,  36694,  36802,  36911,
    37076,  37326,  37626,  37935,  38199,  38397,  38558,  38706,
    38878,  39065,  39266,  39471,  39681,  39899,  40126,  40350,
    40558,  40729,  40881,  41032,  41220,  41447,  41704,  41968,
    42225,  42528,  42870,  43124,  43154,  42798,  42172,  41553,
    41213,  41279,  41589,  41977,  42284,  42458,  42590,  42719,
    42897,  43140,  43427,  43714,  43967,  44171,  44349,  44507,
    44642,  44722,  44758,  44817,  44962,  45229,  45585,  45960,
    46299,  46603,  46899,  47153,  47340,  47400,  47370,  47340,
    47403,  47597,  47877,  48177,  48444,  48668,  48882,  49073,
    49235,  49340,  49403,  49465,  49574,  49742,  49946,  50167,
    50388,  50605,  50829,  51056,  51274,  51475,  51669,  51863,
    52064,  52288,  52529,  52753,  52931,  53036,  53095,  53145,
    53221,  53323,  53441,  53576,  53741,  53939,  54169,  54410,
    54647,  54874,  55102,  55329,  55553,  55774,  55998,  56212,
    56406,  56571,  56712,  56851,  57002,  57160,  57322,  57493,
    57674,  57869,  58076,  58287,  58488,  58672,  58847,  59022,
    59206,  59394,  59588,  59786,  59987,  60188,  60395,  60606,
    60817,  61041,  61275,  61496,  61677,  61785,  61848,  61914,
    62033,  62217,  62448,  62701,  62971,  63274,  63614,  63933,
    64180,  64342,  64447,  64500,  64510,  64434,  64292,  64147,
    64085,  64114,  64200,  64329,  64490,  64694,  64948,  65208,
    65439,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
	 
	 
	 
	// 2 resid 6581
      724,    724,    724,    724,    724,    724,    724,    724,
      724,    728,    728,    728,    728,    728,    728,    728,
      728,    731,    731,    731,    731,    731,    731,    731,
      731,    734,    734,    734,    734,    734,    734,    734,
      737,    737,    737,    737,    737,    737,    737,    741,
      741,    741,    741,    741,    741,    744,    744,    744,
      744,    744,    747,    747,    747,    747,    747,    751,
      751,    751,    751,    751,    754,    754,    754,    754,
      757,    757,    757,    757,    757,    760,    760,    760,
      760,    764,    764,    764,    764,    764,    767,    767,
      767,    767,    770,    770,    770,    770,    770,    774,
      774,    774,    774,    777,    777,    777,    777,    780,
      780,    780,    784,    784,    784,    784,    787,    787,
      787,    790,    790,    790,    793,    793,    793,    797,
      797,    800,    800,    800,    803,    803,    807,    807,
      807,    810,    810,    813,    813,    816,    816,    820,
      823,    823,    826,    826,    830,    830,    833,    833,
      836,    836,    840,    840,    843,    846,    846,    849,
      849,    853,    853,    856,    859,    859,    863,    863,
      866,    869,    869,    872,    876,    876,    879,    882,
      882,    886,    889,    889,    892,    896,    899,    899,
      902,    905,    909,    912,    915,    919,    919,    922,
      925,    928,    932,    935,    938,    942,    945,    952,
      955,    958,    961,    965,    968,    975,    978,    981,
      988,    991,    994,    998,   1004,   1008,   1011,   1014,
     1021,   1024,   1027,   1031,   1034,   1037,   1044,   1047,
     1050,   1054,   1057,   1064,   1067,   1070,   1073,   1080,
     1083,   1087,   1090,   1096,   1100,   1106,   1110,   1116,
     1120,   1126,   1129,   1136,   1143,   1146,   1152,   1159,
     1166,   1172,   1179,   1185,   1192,   1199,   1205,   1215,
     1222,   1228,   1238,   1245,   1255,   1264,   1274,   1284,
     1294,   1304,   1314,   1324,   1334,   1347,   1357,   1370,
     1383,   1393,   1406,   1419,   1432,   1442,   1456,   1469,
     1482,   1495,   1508,   1521,   1535,   1548,   1561,   1574,
     1587,   1600,   1614,   1630,   1643,   1656,   1673,   1686,
     1703,   1716,   1732,   1749,   1765,   1782,   1798,   1815,
     1831,   1848,   1864,   1884,   1900,   1920,   1940,   1956,
     1976,   1996,   2016,   2039,   2058,   2078,   2101,   2124,
     2147,   2167,   2193,   2216,   2240,   2266,   2289,   2315,
     2342,   2368,   2394,   2421,   2450,   2480,   2506,   2536,
     2569,   2599,   2628,   2661,   2691,   2724,   2757,   2790,
     2823,   2859,   2892,   2928,   2961,   2997,   3033,   3070,
     3106,   3142,   3182,   3218,   3257,   3297,   3333,   3373,
     3412,   3452,   3495,   3534,   3577,   3617,   3659,   3702,
     3745,   3788,   3831,   3873,   3916,   3962,   4005,   4051,
     4094,   4140,   4186,   4233,   4279,   4325,   4374,   4420,
     4470,   4516,   4565,   4611,   4661,   4710,   4760,   4809,
     4858,   4911,   4961,   5010,   5063,   5112,   5165,   5218,
     5270,   5323,   5376,   5432,   5491,   5550,   5613,   5675,
     5741,   5807,   5873,   5942,   6011,   6081,   6153,   6226,
     6301,   6377,   6453,   6529,   6604,   6683,   6762,   6842,
     6921,   7003,   7082,   7164,   7247,   7329,   7411,   7494,
     7576,   7659,   7741,   7823,   7909,   7995,   8080,   8166,
     8255,   8340,   8429,   8518,   8611,   8699,   8792,   8881,
     8976,   9068,   9161,   9256,   9352,   9447,   9543,   9638,
     9737,   9836,   9935,  10034,  10132,  10235,  10333,  10436,
    10541,  10643,  10745,  10851,  10956,  11061,  11170,  11276,
    11384,  11493,  11602,  11710,  11822,  11931,  12043,  12155,
    12270,  12382,  12498,  12613,  12728,  12844,  12959,  13077,
    13196,  13315,  13433,  13552,  13674,  13796,  13917,  14039,
    14165,  14290,  14418,  14550,  14688,  14827,  14968,  15113,
    15262,  15410,  15558,  15710,  15861,  16013,  16164,  16319,
    16470,  16619,  16774,  16928,  17087,  17251,  17423,  17600,
    17788,  17999,  18246,  18510,  18776,  19047,  19327,  19616,
    15153,  15324,  15495,  15660,  15812,  15953,  16092,  16230,
    16368,  16503,  16638,  16774,  16909,  17044,  17179,  17317,
    17459,  17600,  17742,  17887,  18035,  18180,  18328,  18477,
    18625,  18773,  18918,  19063,  19208,  19350,  19491,  19626,
    19765,  19896,  20025,  20153,  20282,  20404,  20529,  20651,
    20773,  20891,  21013,  21132,  21254,  21372,  21494,  21616,
    21741,  21863,  21988,  22113,  22235,  22361,  22486,  22611,
    22736,  22861,  22983,  23108,  23230,  23352,  23474,  23596,
    23718,  23836,  23955,  24074,  24192,  24311,  24429,  24548,
    24666,  24782,  24900,  25019,  25134,  25253,  25371,  25487,
    25605,  25721,  25839,  25954,  26070,  26188,  26304,  26422,
    26538,  26656,  26771,  26887,  27005,  27121,  27239,  27355,
    27473,  27588,  27704,  27822,  27941,  28056,  28175,  28290,
    28409,  28527,  28646,  28761,  28880,  28998,  29117,  29236,
    29354,  29476,  29595,  29713,  29832,  29954,  30072,  30194,
    30316,  30435,  30556,  30678,  30800,  30922,  31047,  31169,
    31294,  31416,  31541,  31663,  31789,  31914,  32039,  32164,
    32289,  32418,  32543,  32668,  32797,  32922,  33050,  33179,
    33304,  33432,  33561,  33689,  33818,  33946,  34075,  34203,
    34332,  34463,  34592,  34720,  34849,  34981,  35109,  35241,
    35369,  35498,  35630,  35758,  35890,  36022,  36150,  36282,
    36410,  36542,  36671,  36802,  36934,  37063,  37194,  37323,
    37455,  37583,  37715,  37843,  37975,  38103,  38235,  38364,
    38496,  38624,  38752,  38884,  39013,  39141,  39270,  39398,
    39530,  39658,  39787,  39919,  40050,  40182,  40314,  40446,
    40581,  40716,  40848,  40983,  41121,  41256,  41391,  41526,
    41665,  41800,  41938,  42076,  42211,  42350,  42488,  42623,
    42761,  42900,  43035,  43173,  43308,  43443,  43582,  43717,
    43852,  43987,  44122,  44254,  44389,  44521,  44652,  44784,
    44916,  45048,  45176,  45305,  45433,  45562,  45687,  45812,
    45937,  46059,  46181,  46303,  46425,  46543,  46659,  46777,
    46892,  47004,  47120,  47228,  47340,  47449,  47555,  47660,
    47765,  47868,  47966,  48068,  48164,  48263,  48358,  48454,
    48549,  48642,  48734,  48823,  48912,  49001,  49090,  49175,
    49261,  49347,  49429,  49515,  49597,  49676,  49758,  49837,
    49916,  49996,  50071,  50147,  50223,  50299,  50374,  50450,
    50523,  50595,  50668,  50740,  50813,  50882,  50954,  51023,
    51093,  51162,  51231,  51300,  51369,  51438,  51504,  51573,
    51639,  51705,  51774,  51840,  51906,  51972,  52041,  52107,
    52173,  52239,  52305,  52371,  52440,  52506,  52572,  52638,
    52707,  52773,  52838,  52904,  52970,  53036,  53102,  53168,
    53234,  53296,  53362,  53425,  53491,  53553,  53616,  53678,
    53741,  53804,  53866,  53929,  53991,  54051,  54113,  54173,
    54232,  54291,  54354,  54410,  54469,  54528,  54588,  54644,
    54703,  54759,  54815,  54871,  54927,  54983,  55039,  55095,
    55148,  55204,  55256,  55309,  55362,  55415,  55467,  55517,
    55569,  55619,  55671,  55721,  55770,  55820,  55869,  55915,
    55965,  56011,  56057,  56103,  56149,  56195,  56241,  56284,
    56330,  56373,  56416,  56459,  56498,  56541,  56581,  56620,
    56660,  56699,  56739,  56778,  56815,  56851,  56890,  56927,
    56963,  56996,  57032,  57068,  57101,  57134,  57167,  57200,
    57233,  57266,  57299,  57328,  57361,  57391,  57421,  57450,
    57480,  57510,  57539,  57569,  57595,  57625,  57651,  57681,
    57707,  57734,  57763,  57790,  57816,  57842,  57869,  57892,
    57918,  57944,  57968,  57994,  58017,  58043,  58066,  58093,
    58116,  58139,  58165,  58188,  58211,  58234,  58257,  58280,
    58307,  58330,  58350,  58373,  58396,  58416,  58439,  58458,
    58481,  58501,  58521,  58541,  58560,  58580,  58597,  58616,
    58636,  58653,  58669,  58689,  58705,  58722,  58738,  58755,
    58771,  58788,  58804,  58821,  58834,  58850,  58864,  58880,
    58893,  58910,  58923,  58936,  58952,  58966,  58979,  58992,
    59005,  59018,  59032,  59045,  59058,  59071,  59084,  59097,
    59107,  59120,  59134,  59144,  59157,  59170,  59180,  59193,
    59206,  59216,  59229,  59239,  59252,  59265,  59275,  59288,
	 
	 

	// 3 resid 6581/2
      362,    362,    362,    362,    362,    362,    362,    362,
      362,    364,    364,    364,    364,    364,    364,    364,
      364,    365,    365,    365,    365,    365,    365,    365,
      365,    367,    367,    367,    367,    367,    367,    367,
      368,    368,    368,    368,    368,    368,    368,    370,
      370,    370,    370,    370,    370,    372,    372,    372,
      372,    372,    373,    373,    373,    373,    373,    375,
      375,    375,    375,    375,    377,    377,    377,    377,
      378,    378,    378,    378,    378,    380,    380,    380,
      380,    382,    382,    382,    382,    382,    383,    383,
      383,    383,    385,    385,    385,    385,    385,    387,
      387,    387,    387,    388,    388,    388,    388,    390,
      390,    390,    392,    392,    392,    392,    393,    393,
      393,    395,    395,    395,    396,    396,    396,    398,
      398,    400,    400,    400,    401,    401,    403,    403,
      403,    405,    405,    406,    406,    408,    408,    410,
      411,    411,    413,    413,    415,    415,    416,    416,
      418,    418,    420,    420,    421,    423,    423,    424,
      424,    426,    426,    428,    429,    429,    431,    431,
      433,    434,    434,    436,    438,    438,    439,    441,
      441,    443,    444,    444,    446,    448,    449,    449,
      451,    452,    454,    456,    457,    459,    459,    461,
      462,    464,    466,    467,    469,    471,    472,    476,
      477,    479,    480,    482,    484,    487,    489,    490,
      494,    495,    497,    499,    502,    504,    505,    507,
      510,    512,    513,    515,    517,    518,    522,    523,
      525,    527,    528,    532,    533,    535,    536,    540,
      541,    543,    545,    548,    550,    553,    555,    558,
      560,    563,    564,    568,    571,    573,    576,    579,
      583,    586,    589,    592,    596,    599,    602,    607,
      611,    614,    619,    622,    627,    632,    637,    642,
      647,    652,    657,    662,    667,    673,    678,    685,
      691,    696,    703,    709,    716,    721,    728,    734,
      741,    747,    754,    760,    767,    774,    780,    787,
      793,    800,    807,    815,    821,    828,    836,    843,
      851,    858,    866,    874,    882,    891,    899,    907,
      915,    924,    932,    942,    950,    960,    970,    978,
      988,    998,   1008,   1019,   1029,   1039,   1050,   1062,
     1073,   1083,   1096,   1108,   1120,   1133,   1144,   1157,
     1171,   1184,   1197,   1210,   1225,   1240,   1253,   1268,
     1284,   1299,   1314,   1330,   1345,   1362,   1378,   1395,
     1411,   1429,   1446,   1464,   1480,   1498,   1516,   1535,
     1553,   1571,   1591,   1609,   1628,   1648,   1666,   1686,
     1706,   1726,   1747,   1767,   1788,   1808,   1829,   1851,
     1872,   1894,   1915,   1936,   1958,   1981,   2002,   2025,
     2047,   2070,   2093,   2116,   2139,   2162,   2187,   2210,
     2235,   2258,   2282,   2305,   2330,   2355,   2380,   2404,
     2429,   2455,   2480,   2505,   2531,   2556,   2582,   2609,
     2635,   2661,   2688,   2716,   2745,   2775,   2806,   2837,
     2870,   2903,   2936,   2971,   3005,   3040,   3076,   3113,
     3150,   3188,   3226,   3264,   3302,   3341,   3381,   3421,
     3460,   3501,   3541,   3582,   3623,   3664,   3705,   3747,
     3788,   3829,   3870,   3911,   3954,   3997,   4040,   4083,
     4127,   4170,   4214,   4259,   4305,   4349,   4396,   4440,
     4488,   4534,   4580,   4628,   4676,   4723,   4771,   4819,
     4868,   4918,   4967,   5017,   5066,   5117,   5166,   5218,
     5270,   5321,   5372,   5425,   5478,   5530,   5585,   5638,
     5692,   5746,   5801,   5855,   5911,   5965,   6021,   6077,
     6135,   6191,   6249,   6306,   6364,   6422,   6479,   6538,
     6598,   6657,   6716,   6776,   6837,   6898,   6958,   7019,
     7082,   7145,   7209,   7275,   7344,   7413,   7484,   7556,
     7631,   7705,   7779,   7855,   7930,   8006,   8082,   8159,
     8235,   8309,   8387,   8464,   8543,   8625,   8711,   8800,
     8894,   8999,   9123,   9255,   9388,   9523,   9663,   9808,
     7576,   7662,   7747,   7830,   7906,   7976,   8046,   8115,
     8184,   8251,   8319,   8387,   8454,   8522,   8589,   8658,
     8729,   8800,   8871,   8943,   9017,   9090,   9164,   9238,
     9312,   9386,   9459,   9531,   9604,   9675,   9745,   9813,
     9882,   9948,  10012,  10076,  10141,  10202,  10264,  10325,
    10386,  10445,  10506,  10566,  10627,  10686,  10747,  10808,
    10870,  10931,  10994,  11056,  11117,  11180,  11243,  11305,
    11368,  11430,  11491,  11554,  11615,  11676,  11737,  11798,
    11859,  11918,  11977,  12037,  12096,  12155,  12214,  12274,
    12333,  12391,  12450,  12509,  12567,  12626,  12685,  12743,
    12802,  12860,  12919,  12977,  13035,  13094,  13152,  13211,
    13269,  13328,  13385,  13443,  13502,  13560,  13619,  13677,
    13736,  13794,  13852,  13911,  13970,  14028,  14087,  14145,
    14204,  14263,  14323,  14380,  14440,  14499,  14558,  14618,
    14677,  14738,  14797,  14856,  14916,  14977,  15036,  15097,
    15158,  15217,  15278,  15339,  15400,  15461,  15523,  15584,
    15647,  15708,  15770,  15831,  15894,  15957,  16019,  16082,
    16144,  16209,  16271,  16334,  16398,  16461,  16525,  16589,
    16652,  16716,  16780,  16844,  16909,  16973,  17037,  17101,
    17166,  17231,  17296,  17360,  17424,  17490,  17554,  17620,
    17684,  17749,  17815,  17879,  17945,  18011,  18075,  18141,
    18205,  18271,  18335,  18401,  18467,  18531,  18597,  18661,
    18727,  18791,  18857,  18921,  18987,  19051,  19117,  19182,
    19248,  19312,  19376,  19442,  19506,  19570,  19635,  19699,
    19765,  19829,  19893,  19959,  20025,  20091,  20157,  20223,
    20290,  20358,  20424,  20491,  20560,  20628,  20695,  20763,
    20832,  20900,  20969,  21038,  21105,  21175,  21244,  21311,
    21380,  21450,  21517,  21586,  21654,  21721,  21791,  21858,
    21926,  21993,  22061,  22127,  22194,  22260,  22326,  22392,
    22458,  22524,  22588,  22652,  22716,  22781,  22843,  22906,
    22968,  23029,  23090,  23151,  23212,  23271,  23329,  23388,
    23446,  23502,  23560,  23614,  23670,  23724,  23777,  23830,
    23882,  23934,  23983,  24034,  24082,  24131,  24179,  24227,
    24274,  24321,  24367,  24411,  24456,  24500,  24545,  24587,
    24630,  24673,  24714,  24757,  24798,  24838,  24879,  24918,
    24958,  24998,  25035,  25073,  25111,  25149,  25187,  25225,
    25261,  25297,  25334,  25370,  25406,  25441,  25477,  25511,
    25546,  25581,  25615,  25650,  25684,  25719,  25752,  25786,
    25819,  25852,  25887,  25920,  25953,  25986,  26020,  26053,
    26086,  26119,  26152,  26185,  26220,  26253,  26286,  26319,
    26353,  26386,  26419,  26452,  26485,  26518,  26551,  26584,
    26617,  26648,  26681,  26712,  26745,  26776,  26808,  26839,
    26870,  26902,  26933,  26964,  26995,  27025,  27056,  27086,
    27116,  27145,  27177,  27205,  27234,  27264,  27294,  27322,
    27351,  27379,  27407,  27435,  27463,  27491,  27519,  27547,
    27574,  27602,  27628,  27654,  27681,  27707,  27733,  27758,
    27784,  27809,  27835,  27860,  27885,  27910,  27934,  27957,
    27982,  28005,  28028,  28051,  28074,  28097,  28120,  28142,
    28165,  28186,  28208,  28229,  28249,  28270,  28290,  28310,
    28330,  28349,  28369,  28389,  28407,  28425,  28445,  28463,
    28481,  28498,  28516,  28534,  28550,  28567,  28583,  28600,
    28616,  28633,  28649,  28664,  28680,  28695,  28710,  28725,
    28740,  28755,  28769,  28784,  28797,  28812,  28825,  28840,
    28853,  28867,  28881,  28895,  28908,  28921,  28934,  28946,
    28959,  28972,  28984,  28997,  29008,  29021,  29033,  29046,
    29058,  29069,  29082,  29094,  29105,  29117,  29128,  29140,
    29153,  29165,  29175,  29186,  29198,  29208,  29219,  29229,
    29240,  29250,  29260,  29270,  29280,  29290,  29298,  29308,
    29318,  29326,  29334,  29344,  29352,  29361,  29369,  29377,
    29385,  29394,  29402,  29410,  29417,  29425,  29432,  29440,
    29446,  29455,  29461,  29468,  29476,  29483,  29489,  29496,
    29502,  29509,  29516,  29522,  29529,  29535,  29542,  29548,
    29553,  29560,  29567,  29572,  29578,  29585,  29590,  29596,
    29603,  29608,  29614,  29619,  29626,  29632,  29637,  29644
};

endmodule
