-------------------------------------------------------------------------------
--
-- (C) COPYRIGHT 2010 Gideon's Logic Architectures'
--
-------------------------------------------------------------------------------
-- 
-- Author: Gideon Zweijtzer (gideon.zweijtzer (at) gmail.com)
--
-- Note that this file is copyrighted, and is not supposed to be used in other
-- projects without written permission from the author.
--
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.my_math_pkg.all;

entity sid_filter is
port (
    clock       : in  std_logic;
    reset       : in  std_logic;
    enable      : in  std_logic;

    cfg         : in  unsigned(2 downto 0);
    
    filt_co     : in  unsigned(10 downto 0);
    filt_res    : in  unsigned(3 downto 0);

    valid_in    : in  std_logic := '0';
    error_out   : out std_logic;     
    input       : in  signed(17 downto 0);
    high_pass   : out signed(17 downto 0);
    band_pass   : out signed(17 downto 0);
    low_pass    : out signed(17 downto 0);
	 
    valid_out   : out std_logic;

	 ld_clk      : in  std_logic;
	 ld_addr     : in  std_logic_vector(11 downto 0);
	 ld_data     : in  std_logic_vector(15 downto 0);
	 ld_wr       : in  std_logic
);
end entity;

architecture dsvf of sid_filter is
    type t_word_array is array(0 to (8*1024)-1) of signed(15 downto 0);
    signal coef : t_word_array := 
    (
      -- Config 0
      x"0320", x"0321", x"0322", x"0322", x"0323", x"0323", x"0324", x"0324", x"0325", x"0326", x"0326", x"0327", x"0327", x"0328", x"0328", x"0329",
      x"032A", x"032A", x"032B", x"032B", x"032C", x"032C", x"032D", x"032E", x"032E", x"032F", x"032F", x"0330", x"0330", x"0331", x"0332", x"0332",
      x"0333", x"0333", x"0334", x"0334", x"0335", x"0336", x"0336", x"0337", x"0337", x"0338", x"0338", x"0339", x"033A", x"033A", x"033B", x"033B",
      x"033C", x"033C", x"033D", x"033E", x"033E", x"033F", x"033F", x"0340", x"0340", x"0341", x"0341", x"0342", x"0343", x"0343", x"0344", x"0344",
      x"0345", x"0346", x"0347", x"0348", x"0349", x"034B", x"034C", x"034D", x"034E", x"034F", x"0350", x"0351", x"0353", x"0354", x"0355", x"0356",
      x"0357", x"0358", x"0359", x"035B", x"035C", x"035D", x"035E", x"035F", x"0360", x"0361", x"0362", x"0364", x"0365", x"0366", x"0367", x"0368",
      x"0369", x"036A", x"036C", x"036D", x"036E", x"036F", x"0370", x"0371", x"0372", x"0374", x"0375", x"0376", x"0377", x"0378", x"0379", x"037A",
      x"037C", x"037D", x"037E", x"037F", x"0380", x"0381", x"0382", x"0383", x"0385", x"0386", x"0387", x"0388", x"0389", x"038A", x"038B", x"038D",
      x"038E", x"0391", x"0393", x"0396", x"0399", x"039C", x"039F", x"03A2", x"03A4", x"03A7", x"03AA", x"03AD", x"03B0", x"03B3", x"03B6", x"03B8",
      x"03BB", x"03BE", x"03C1", x"03C4", x"03C7", x"03C9", x"03CC", x"03CF", x"03D2", x"03D5", x"03D8", x"03DB", x"03DD", x"03E0", x"03E3", x"03E6",
      x"03E9", x"03EC", x"03EE", x"03F1", x"03F4", x"03F7", x"03FA", x"03FD", x"03FF", x"0402", x"0405", x"0408", x"040B", x"040E", x"0411", x"0413",
      x"0416", x"0419", x"041C", x"041F", x"0422", x"0424", x"0427", x"042A", x"042D", x"0430", x"0433", x"0436", x"0438", x"043B", x"043E", x"0441",
      x"0444", x"044B", x"0451", x"0458", x"045F", x"0466", x"046D", x"0474", x"047A", x"0481", x"0488", x"048F", x"0496", x"049D", x"04A3", x"04AA",
      x"04B1", x"04B8", x"04BF", x"04C5", x"04CC", x"04D3", x"04DA", x"04E1", x"04E8", x"04EE", x"04F5", x"04FC", x"0503", x"050A", x"0511", x"0517",
      x"051E", x"0525", x"052C", x"0533", x"053A", x"0540", x"0547", x"054E", x"0555", x"055C", x"0562", x"0569", x"0570", x"0577", x"057E", x"0585",
      x"058B", x"0592", x"0599", x"05A0", x"05A7", x"05AE", x"05B4", x"05BB", x"05C2", x"05C9", x"05D0", x"05D7", x"05DD", x"05E4", x"05EB", x"05F2",
      x"05F9", x"060D", x"0622", x"0636", x"064B", x"065F", x"0674", x"0688", x"069D", x"06B1", x"06C5", x"06DA", x"06EE", x"0703", x"0717", x"072C",
      x"0740", x"0755", x"0769", x"077E", x"0792", x"07A7", x"07BB", x"07D0", x"07E4", x"07F9", x"080D", x"0822", x"0836", x"084B", x"085F", x"0874",
      x"0888", x"089C", x"08B1", x"08C5", x"08DA", x"08EE", x"0903", x"0917", x"092C", x"0940", x"0955", x"0969", x"097E", x"0992", x"09A7", x"09BB",
      x"09D0", x"09E4", x"09F9", x"0A0D", x"0A22", x"0A36", x"0A4B", x"0A5F", x"0A74", x"0A88", x"0A9C", x"0AB1", x"0AC5", x"0ADA", x"0AEE", x"0B03",
      x"0B17", x"0B46", x"0B75", x"0BA3", x"0BD2", x"0C01", x"0C2F", x"0C5E", x"0C8D", x"0CBB", x"0CEA", x"0D19", x"0D47", x"0D76", x"0DA4", x"0DD3",
      x"0E02", x"0E30", x"0E5F", x"0E8E", x"0EBC", x"0EEB", x"0F1A", x"0F48", x"0F77", x"0FA6", x"0FD4", x"1003", x"1032", x"1060", x"108F", x"10BD",
      x"10EC", x"111B", x"1149", x"1178", x"11A7", x"11D5", x"1204", x"1233", x"1261", x"1290", x"12BF", x"12ED", x"131C", x"134B", x"1379", x"13A8",
      x"13D7", x"1405", x"1434", x"1462", x"1491", x"14C0", x"14EE", x"151D", x"154C", x"157A", x"15A9", x"15D8", x"1606", x"1635", x"1664", x"1692",
      x"16C1", x"1711", x"1760", x"17B0", x"17FF", x"184F", x"189F", x"18EE", x"193E", x"198E", x"19DD", x"1A2D", x"1A7D", x"1ACC", x"1B1C", x"1B6C",
      x"1BBB", x"1C0B", x"1C5A", x"1CAA", x"1CFA", x"1D49", x"1D99", x"1DE9", x"1E38", x"1E88", x"1ED8", x"1F27", x"1F77", x"1FC7", x"2016", x"2066",
      x"20B5", x"211C", x"2182", x"21E9", x"224F", x"22B5", x"231C", x"2382", x"23E9", x"244F", x"24B5", x"251C", x"2582", x"25E9", x"264F", x"26B5",
      x"271C", x"2782", x"27E9", x"284F", x"28B5", x"291C", x"2982", x"29E9", x"2A4F", x"2AB5", x"2B1C", x"2B82", x"2BE9", x"2C4F", x"2CB5", x"2D1C",
      x"2D82", x"2DFF", x"2E7D", x"2EFA", x"2F77", x"2FF4", x"3071", x"30EE", x"316B", x"31E9", x"3266", x"32E3", x"3360", x"33DD", x"345A", x"34D8",
      x"3555", x"35D2", x"364F", x"36CC", x"3749", x"37C7", x"3844", x"38C1", x"393E", x"39BB", x"3A38", x"3AB5", x"3B33", x"3BB0", x"3C2D", x"3CAA",
      x"3D27", x"3DC6", x"3E66", x"3F05", x"3FA4", x"4044", x"40E3", x"4182", x"4222", x"42C1", x"4360", x"43FF", x"449F", x"453E", x"45DD", x"467D",
      x"471C", x"47D2", x"4888", x"493E", x"49F4", x"4AAA", x"4B60", x"4C16", x"4CCC", x"4DDD", x"4EEE", x"4FFF", x"5110", x"5248", x"5381", x"54B9",
      x"416B", x"4222", x"42D8", x"438E", x"4444", x"44DB", x"4573", x"460B", x"46A2", x"473A", x"47D2", x"486A", x"4901", x"4999", x"4A31", x"4AC8",
      x"4B60", x"4BFF", x"4C9F", x"4D3E", x"4DDD", x"4E7D", x"4F1C", x"4FBB", x"505A", x"50FA", x"5199", x"5238", x"52D8", x"5377", x"5416", x"54B5",
      x"5555", x"55DD", x"5666", x"56EE", x"5777", x"57FF", x"5888", x"5910", x"5999", x"5A21", x"5AAA", x"5B33", x"5BBB", x"5C44", x"5CCC", x"5D55",
      x"5DDD", x"5E66", x"5EEE", x"5F77", x"5FFF", x"6088", x"6110", x"6199", x"6221", x"62AA", x"6333", x"63BB", x"6444", x"64CC", x"6555", x"65DD",
      x"6666", x"66E9", x"676B", x"67EE", x"6871", x"68F4", x"6977", x"69FA", x"6A7C", x"6AFF", x"6B82", x"6C05", x"6C88", x"6D0B", x"6D8E", x"6E10",
      x"6E93", x"6F16", x"6F99", x"701C", x"709F", x"7121", x"71A4", x"7227", x"72AA", x"732D", x"73B0", x"7432", x"74B5", x"7538", x"75BB", x"763E",
      x"76C1", x"7744", x"77C6", x"7849", x"78CC", x"794F", x"79D2", x"7A55", x"7AD7", x"7B5A", x"7BDD", x"7C60", x"7CE3", x"7D66", x"7DE8", x"7E6B",
      x"7EEE", x"7F71", x"7FF4", x"8077", x"80FA", x"817C", x"81FF", x"8282", x"8305", x"8388", x"840B", x"848D", x"8510", x"8593", x"8616", x"8699",
      x"871C", x"87AA", x"8838", x"88C6", x"8955", x"89E3", x"8A71", x"8AFF", x"8B8D", x"8C1C", x"8CAA", x"8D38", x"8DC6", x"8E55", x"8EE3", x"8F71",
      x"8FFF", x"908D", x"911C", x"91AA", x"9238", x"92C6", x"9355", x"93E3", x"9471", x"94FF", x"958D", x"961C", x"96AA", x"9738", x"97C6", x"9855",
      x"98E3", x"9971", x"99FF", x"9A8D", x"9B1C", x"9BAA", x"9C38", x"9CC6", x"9D55", x"9DE3", x"9E71", x"9EFF", x"9F8D", x"A01C", x"A0AA", x"A138",
      x"A1C6", x"A255", x"A2E3", x"A371", x"A3FF", x"A48D", x"A51C", x"A5AA", x"A638", x"A6C6", x"A755", x"A7E3", x"A871", x"A8FF", x"A98D", x"AA1C",
      x"AAAA", x"AB38", x"ABC6", x"AC54", x"ACE3", x"AD71", x"ADFF", x"AE8D", x"AF1C", x"AFAA", x"B038", x"B0C6", x"B154", x"B1E3", x"B271", x"B2FF",
      x"B38D", x"B41C", x"B4AA", x"B538", x"B5C6", x"B654", x"B6E3", x"B771", x"B7FF", x"B88D", x"B91C", x"B9AA", x"BA38", x"BAC6", x"BB54", x"BBE3",
      x"BC71", x"BCFF", x"BD8D", x"BE1C", x"BEAA", x"BF38", x"BFC6", x"C054", x"C0E3", x"C171", x"C1FF", x"C28D", x"C31C", x"C3AA", x"C438", x"C4C6",
      x"C554", x"C5E3", x"C671", x"C6FF", x"C78D", x"C81C", x"C8AA", x"C938", x"C9C6", x"CA54", x"CAE3", x"CB71", x"CBFF", x"CC8D", x"CD1C", x"CDAA",
      x"CE38", x"CE8D", x"CEE3", x"CF38", x"CF8D", x"CFE3", x"D038", x"D08D", x"D0E3", x"D138", x"D18D", x"D1E3", x"D238", x"D28D", x"D2E3", x"D338",
      x"D38D", x"D3E3", x"D438", x"D48D", x"D4E3", x"D538", x"D58D", x"D5E3", x"D638", x"D68D", x"D6E3", x"D738", x"D78D", x"D7E3", x"D838", x"D88D",
      x"D8E3", x"D938", x"D98D", x"D9E3", x"DA38", x"DA8D", x"DAE3", x"DB38", x"DB8D", x"DBE3", x"DC38", x"DC8D", x"DCE3", x"DD38", x"DD8D", x"DDE3",
      x"DE38", x"DE8D", x"DEE3", x"DF38", x"DF8D", x"DFE3", x"E038", x"E08D", x"E0E3", x"E138", x"E18D", x"E1E3", x"E238", x"E28D", x"E2E3", x"E338",
      x"E38D", x"E3CC", x"E40A", x"E449", x"E488", x"E4C6", x"E505", x"E543", x"E582", x"E5C0", x"E5FF", x"E63E", x"E67C", x"E6BB", x"E6F9", x"E738",
      x"E777", x"E7B5", x"E7F4", x"E832", x"E871", x"E8AF", x"E8EE", x"E92D", x"E96B", x"E9AA", x"E9E8", x"EA27", x"EA65", x"EAA4", x"EAE3", x"EB21",
      x"EB60", x"EB9E", x"EBDD", x"EC1B", x"EC5A", x"EC99", x"ECD7", x"ED16", x"ED54", x"ED93", x"EDD2", x"EE10", x"EE4F", x"EE8D", x"EECC", x"EF0A",
      x"EF49", x"EF88", x"EFC6", x"F005", x"F043", x"F082", x"F0C0", x"F0FF", x"F13E", x"F17C", x"F1BB", x"F1F9", x"F238", x"F276", x"F2B5", x"F2F4",
      x"F332", x"F354", x"F376", x"F399", x"F3BB", x"F3DD", x"F3FF", x"F421", x"F443", x"F465", x"F488", x"F4AA", x"F4CC", x"F4EE", x"F510", x"F532",
      x"F554", x"F576", x"F599", x"F5BB", x"F5DD", x"F5FF", x"F621", x"F643", x"F665", x"F688", x"F6AA", x"F6CC", x"F6EE", x"F710", x"F732", x"F754",
      x"F776", x"F799", x"F7BB", x"F7DD", x"F7FF", x"F821", x"F843", x"F865", x"F888", x"F8AA", x"F8CC", x"F8EE", x"F910", x"F932", x"F954", x"F976",
      x"F999", x"F9BB", x"F9DD", x"F9FF", x"FA21", x"FA43", x"FA65", x"FA88", x"FAAA", x"FACC", x"FAEE", x"FB10", x"FB32", x"FB54", x"FB76", x"FB99",
      x"FBBB", x"FBCC", x"FBDD", x"FBEE", x"FC00", x"FC11", x"FC22", x"FC33", x"FC44", x"FC56", x"FC67", x"FC78", x"FC89", x"FC9A", x"FCAC", x"FCBD",
      x"FCCE", x"FCDF", x"FCF0", x"FD02", x"FD13", x"FD24", x"FD35", x"FD46", x"FD58", x"FD69", x"FD7A", x"FD8B", x"FD9C", x"FDAE", x"FDBF", x"FDD0",
      x"FDE1", x"FDF2", x"FE04", x"FE15", x"FE26", x"FE37", x"FE48", x"FE5A", x"FE6B", x"FE7C", x"FE8D", x"FE9E", x"FEB0", x"FEC1", x"FED2", x"FEE3",
      x"FEF4", x"FF06", x"FF17", x"FF28", x"FF39", x"FF4A", x"FF5C", x"FF6D", x"FF7E", x"FF8F", x"FFA0", x"FFB2", x"FFC3", x"FFD4", x"FFE5", x"FFF6",

      -- Config 1
      x"0005", x"000A", x"000F", x"0013", x"0018", x"001D", x"0023", x"0028", x"002D", x"0032", x"0036", x"003B", x"0040", x"0046", x"004B", x"0050",
      x"0055", x"0059", x"005E", x"0063", x"0069", x"006E", x"0073", x"0078", x"007C", x"0081", x"0086", x"008C", x"0091", x"0096", x"009B", x"009F",
      x"00A4", x"00A9", x"00AF", x"00B4", x"00B9", x"00BE", x"00C2", x"00C7", x"00CC", x"00D2", x"00D7", x"00DC", x"00E1", x"00E5", x"00EA", x"00EF",
      x"00F5", x"00FA", x"00FF", x"0104", x"0108", x"010D", x"0112", x"0118", x"011D", x"0122", x"0127", x"012B", x"0130", x"0135", x"013B", x"0140",
      x"0145", x"014A", x"014E", x"0153", x"0158", x"015E", x"0163", x"0168", x"016D", x"0171", x"0176", x"017B", x"0181", x"0186", x"018B", x"0190",
      x"0194", x"0199", x"019E", x"01A4", x"01A9", x"01AE", x"01B3", x"01B7", x"01BC", x"01C1", x"01C7", x"01CC", x"01D1", x"01D6", x"01DA", x"01DF",
      x"01E4", x"01EA", x"01EF", x"01F4", x"01F9", x"01FD", x"0202", x"0207", x"020D", x"0212", x"0217", x"021C", x"0220", x"0225", x"022A", x"0230",
      x"0235", x"023A", x"023E", x"0243", x"0248", x"024D", x"0253", x"0258", x"025D", x"0261", x"0266", x"026B", x"0270", x"0276", x"027B", x"0280",
      x"0284", x"0289", x"028E", x"0293", x"0299", x"029E", x"02A3", x"02A7", x"02AC", x"02B1", x"02B6", x"02BC", x"02C1", x"02C6", x"02CA", x"02CF",
      x"02D4", x"02D9", x"02DF", x"02E4", x"02E9", x"02ED", x"02F2", x"02F7", x"02FC", x"0302", x"0307", x"030C", x"0310", x"0315", x"031A", x"031F",
      x"0325", x"032A", x"032F", x"0333", x"0338", x"033D", x"0342", x"0348", x"034D", x"0352", x"0356", x"035B", x"0360", x"0365", x"036B", x"0370",
      x"0375", x"0379", x"037E", x"0383", x"0388", x"038E", x"0393", x"0398", x"039C", x"03A1", x"03A6", x"03AB", x"03B1", x"03B6", x"03BB", x"03BF",
      x"03C4", x"03C9", x"03CE", x"03D4", x"03D9", x"03DE", x"03E2", x"03E7", x"03EC", x"03F1", x"03F7", x"03FC", x"0401", x"0405", x"040A", x"040F",
      x"0414", x"041A", x"041F", x"0424", x"0428", x"042D", x"0432", x"0437", x"043D", x"0442", x"0447", x"044B", x"0450", x"0455", x"045A", x"0460",
      x"0465", x"046A", x"046E", x"0473", x"0478", x"047D", x"0483", x"0488", x"048C", x"0491", x"0496", x"049B", x"04A0", x"04A6", x"04AB", x"04AF",
      x"04B4", x"04B9", x"04BE", x"04C3", x"04C9", x"04CE", x"04D2", x"04D7", x"04DC", x"04E1", x"04E6", x"04EC", x"04F1", x"04F5", x"04FA", x"04FF",
      x"0504", x"0509", x"050F", x"0514", x"0518", x"051D", x"0522", x"0527", x"052C", x"0532", x"0537", x"053B", x"0540", x"0545", x"054A", x"054F",
      x"0555", x"055A", x"055E", x"0563", x"0568", x"056D", x"0572", x"0578", x"057D", x"0581", x"0586", x"058B", x"0590", x"0595", x"059B", x"05A0",
      x"05A4", x"05A9", x"05AE", x"05B3", x"05B8", x"05BE", x"05C3", x"05C7", x"05CC", x"05D1", x"05D6", x"05DB", x"05E1", x"05E5", x"05EA", x"05EF",
      x"05F4", x"05F9", x"05FE", x"0604", x"0608", x"060D", x"0612", x"0617", x"061C", x"0621", x"0627", x"062B", x"0630", x"0635", x"063A", x"063F",
      x"0644", x"064A", x"064E", x"0653", x"0658", x"065D", x"0662", x"0667", x"066D", x"0671", x"0676", x"067B", x"0680", x"0685", x"068A", x"0690",
      x"0694", x"0699", x"069E", x"06A3", x"06A8", x"06AD", x"06B3", x"06B7", x"06BC", x"06C1", x"06C6", x"06CB", x"06D0", x"06D5", x"06DA", x"06DF",
      x"06E4", x"06E9", x"06EE", x"06F3", x"06F8", x"06FD", x"0702", x"0707", x"070C", x"0711", x"0716", x"071B", x"0720", x"0725", x"072A", x"072F",
      x"0734", x"0739", x"073E", x"0743", x"0748", x"074D", x"0752", x"0757", x"075C", x"0761", x"0766", x"076B", x"0770", x"0775", x"077A", x"077F",
      x"0784", x"0789", x"078E", x"0793", x"0798", x"079D", x"07A2", x"07A7", x"07AC", x"07B1", x"07B6", x"07BB", x"07C0", x"07C5", x"07CA", x"07CF",
      x"07D4", x"07D9", x"07DE", x"07E3", x"07E8", x"07ED", x"07F2", x"07F7", x"07FC", x"0801", x"0806", x"080B", x"0810", x"0815", x"081A", x"081F",
      x"0824", x"0829", x"082E", x"0833", x"0838", x"083D", x"0842", x"0847", x"084C", x"0851", x"0856", x"085B", x"0860", x"0865", x"086A", x"086F",
      x"0874", x"0879", x"087E", x"0883", x"0888", x"088D", x"0892", x"0897", x"089C", x"08A1", x"08A6", x"08AB", x"08B0", x"08B5", x"08BA", x"08BF",
      x"08C4", x"08C9", x"08CE", x"08D3", x"08D8", x"08DD", x"08E2", x"08E7", x"08EC", x"08F1", x"08F6", x"08FB", x"0900", x"0905", x"090A", x"090F",
      x"0914", x"0919", x"091E", x"0923", x"0928", x"092D", x"0932", x"0937", x"093C", x"0941", x"0946", x"094B", x"0950", x"0955", x"095A", x"095F",
      x"0964", x"0969", x"096E", x"0973", x"0978", x"097D", x"0982", x"0987", x"098C", x"0991", x"0996", x"099B", x"09A0", x"09A5", x"09AA", x"09AF",
      x"09B4", x"09B9", x"09BE", x"09C3", x"09C8", x"09CD", x"09D2", x"09D7", x"09DC", x"09E1", x"09E6", x"09EB", x"09F0", x"09F5", x"09FA", x"09FF",
      x"0A04", x"0A09", x"0A0E", x"0A13", x"0A18", x"0A1D", x"0A22", x"0A27", x"0A2C", x"0A31", x"0A36", x"0A3B", x"0A40", x"0A45", x"0A4A", x"0A4F",
      x"0A54", x"0A59", x"0A5E", x"0A63", x"0A68", x"0A6D", x"0A72", x"0A77", x"0A7C", x"0A81", x"0A86", x"0A8B", x"0A90", x"0A95", x"0A9A", x"0A9F",
      x"0AA4", x"0AA9", x"0AAE", x"0AB3", x"0AB8", x"0ABD", x"0AC2", x"0AC7", x"0ACC", x"0AD1", x"0AD6", x"0ADB", x"0AE0", x"0AE5", x"0AEA", x"0AEF",
      x"0AF4", x"0AF9", x"0AFE", x"0B03", x"0B08", x"0B0D", x"0B12", x"0B17", x"0B1C", x"0B21", x"0B26", x"0B2B", x"0B30", x"0B35", x"0B3A", x"0B3F",
      x"0B44", x"0B49", x"0B4E", x"0B53", x"0B58", x"0B5D", x"0B62", x"0B67", x"0B6C", x"0B71", x"0B76", x"0B7B", x"0B80", x"0B85", x"0B8A", x"0B8F",
      x"0B94", x"0B99", x"0B9E", x"0BA3", x"0BA8", x"0BAD", x"0BB2", x"0BB7", x"0BBC", x"0BC1", x"0BC6", x"0BCB", x"0BD0", x"0BD5", x"0BDA", x"0BDF",
      x"0BE4", x"0BE9", x"0BEE", x"0BF3", x"0BF8", x"0BFD", x"0C02", x"0C07", x"0C0C", x"0C11", x"0C16", x"0C1B", x"0C20", x"0C25", x"0C2A", x"0C2F",
      x"0C34", x"0C39", x"0C3E", x"0C43", x"0C48", x"0C4D", x"0C52", x"0C57", x"0C5C", x"0C61", x"0C66", x"0C6B", x"0C70", x"0C75", x"0C7A", x"0C7F",
      x"0C84", x"0C89", x"0C8E", x"0C93", x"0C98", x"0C9D", x"0CA2", x"0CA7", x"0CAC", x"0CB1", x"0CB6", x"0CBB", x"0CC0", x"0CC5", x"0CCA", x"0CCF",
      x"0CD4", x"0CD9", x"0CDE", x"0CE3", x"0CE8", x"0CED", x"0CF2", x"0CF7", x"0CFC", x"0D01", x"0D06", x"0D0B", x"0D10", x"0D15", x"0D1A", x"0D1F",
      x"0D24", x"0D29", x"0D2E", x"0D33", x"0D38", x"0D3D", x"0D42", x"0D47", x"0D4C", x"0D51", x"0D56", x"0D5B", x"0D60", x"0D65", x"0D6A", x"0D6F",
      x"0D74", x"0D79", x"0D7E", x"0D83", x"0D88", x"0D8D", x"0D92", x"0D97", x"0D9C", x"0DA1", x"0DA6", x"0DAB", x"0DB0", x"0DB5", x"0DBA", x"0DBF",
      x"0DC4", x"0DC9", x"0DCE", x"0DD3", x"0DD8", x"0DDD", x"0DE2", x"0DE7", x"0DEC", x"0DF1", x"0DF6", x"0DFB", x"0E00", x"0E05", x"0E0A", x"0E0F",
      x"0E14", x"0E19", x"0E1E", x"0E23", x"0E28", x"0E2D", x"0E32", x"0E37", x"0E3C", x"0E41", x"0E46", x"0E4B", x"0E50", x"0E55", x"0E5A", x"0E5F",
      x"0E64", x"0E69", x"0E6E", x"0E73", x"0E78", x"0E7D", x"0E82", x"0E87", x"0E8C", x"0E91", x"0E96", x"0E9B", x"0EA0", x"0EA5", x"0EAA", x"0EAF",
      x"0EB4", x"0EB9", x"0EBE", x"0EC3", x"0EC8", x"0ECD", x"0ED2", x"0ED7", x"0EDC", x"0EE1", x"0EE6", x"0EEB", x"0EF0", x"0EF5", x"0EFA", x"0EFF",
      x"0F04", x"0F09", x"0F0E", x"0F13", x"0F18", x"0F1D", x"0F22", x"0F27", x"0F2C", x"0F31", x"0F36", x"0F3B", x"0F40", x"0F45", x"0F4A", x"0F4F",
      x"0F54", x"0F59", x"0F5E", x"0F63", x"0F68", x"0F6D", x"0F72", x"0F77", x"0F7C", x"0F81", x"0F86", x"0F8B", x"0F90", x"0F95", x"0F9A", x"0F9F",
      x"0FA4", x"0FA9", x"0FAE", x"0FB3", x"0FB8", x"0FBD", x"0FC1", x"0FC7", x"0FCC", x"0FD1", x"0FD6", x"0FDB", x"0FE0", x"0FE4", x"0FEA", x"0FEF",
      x"0FF4", x"0FF9", x"0FFE", x"1002", x"1007", x"100D", x"1012", x"1017", x"101C", x"1020", x"1025", x"102A", x"1030", x"1035", x"103A", x"103F",
      x"1043", x"1048", x"104D", x"1053", x"1058", x"105D", x"1061", x"1066", x"106B", x"1070", x"1076", x"107B", x"107F", x"1084", x"1089", x"108E",
      x"1093", x"1099", x"109D", x"10A2", x"10A7", x"10AC", x"10B1", x"10B6", x"10BC", x"10C0", x"10C5", x"10CA", x"10CF", x"10D4", x"10D9", x"10DE",
      x"10E3", x"10E8", x"10ED", x"10F2", x"10F7", x"10FC", x"1101", x"1106", x"110B", x"1110", x"1115", x"111A", x"111F", x"1124", x"1129", x"112E",
      x"1133", x"1138", x"113D", x"1142", x"1147", x"114C", x"1151", x"1156", x"115B", x"1160", x"1165", x"116A", x"116F", x"1174", x"1179", x"117E",
      x"1183", x"1188", x"118D", x"1192", x"1197", x"119C", x"11A1", x"11A6", x"11AB", x"11B0", x"11B5", x"11BA", x"11BF", x"11C4", x"11C9", x"11CE",
      x"11D3", x"11D8", x"11DD", x"11E2", x"11E7", x"11EC", x"11F1", x"11F6", x"11FB", x"1200", x"1205", x"120A", x"120F", x"1214", x"1219", x"121E",
      x"1223", x"1228", x"122D", x"1232", x"1237", x"123C", x"1241", x"1246", x"124B", x"1250", x"1255", x"125A", x"125F", x"1264", x"1269", x"126E",
      x"1273", x"1278", x"127D", x"1282", x"1287", x"128C", x"1291", x"1296", x"129B", x"12A0", x"12A5", x"12AA", x"12AF", x"12B4", x"12B9", x"12BE",
      x"12C3", x"12C8", x"12CD", x"12D2", x"12D7", x"12DC", x"12E1", x"12E6", x"12EB", x"12F0", x"12F5", x"12FA", x"12FF", x"1304", x"1309", x"130E",
      x"1313", x"1318", x"131D", x"1322", x"1327", x"132C", x"1331", x"1336", x"133B", x"1340", x"1345", x"134A", x"134F", x"1354", x"1359", x"135E",
      x"1363", x"1368", x"136D", x"1372", x"1377", x"137C", x"1381", x"1386", x"138B", x"1390", x"1395", x"139A", x"139F", x"13A4", x"13A9", x"13AE",
      x"13B3", x"13B8", x"13BD", x"13C2", x"13C7", x"13CC", x"13D1", x"13D6", x"13DB", x"13E0", x"13E5", x"13EA", x"13EF", x"13F4", x"13F9", x"13FE",

      -- Config 2
      x"0006", x"000D", x"0013", x"001A", x"0020", x"0027", x"002D", x"0034", x"003A", x"0041", x"0047", x"004E", x"0054", x"005B", x"0062", x"0068",
      x"006F", x"0075", x"007C", x"0082", x"0089", x"008F", x"0096", x"009C", x"00A3", x"00A9", x"00B0", x"00B6", x"00BD", x"00C4", x"00CA", x"00D0",
      x"00D7", x"00DE", x"00E4", x"00EB", x"00F1", x"00F8", x"00FE", x"0105", x"010B", x"0112", x"0118", x"011F", x"0126", x"012C", x"0132", x"0139",
      x"0140", x"0146", x"014D", x"0153", x"015A", x"0160", x"0167", x"016D", x"0174", x"017A", x"0181", x"0187", x"018E", x"0194", x"019B", x"01A2",
      x"01A8", x"01AF", x"01B5", x"01BC", x"01C2", x"01C9", x"01CF", x"01D6", x"01DC", x"01E3", x"01E9", x"01F0", x"01F6", x"01FD", x"0204", x"020A",
      x"0210", x"0217", x"021E", x"0224", x"022B", x"0231", x"0238", x"023E", x"0245", x"024B", x"0252", x"0258", x"025F", x"0266", x"026C", x"0272",
      x"0279", x"0280", x"0286", x"028D", x"0293", x"029A", x"02A0", x"02A7", x"02AD", x"02B4", x"02BA", x"02C1", x"02C7", x"02CE", x"02D4", x"02DB",
      x"02E2", x"02E8", x"02EE", x"02F5", x"02FC", x"0302", x"0309", x"030F", x"0316", x"031C", x"0323", x"0329", x"0330", x"0336", x"033D", x"0344",
      x"034A", x"0350", x"0357", x"035E", x"0364", x"036B", x"0371", x"0378", x"037E", x"0385", x"038B", x"0392", x"0398", x"039F", x"03A5", x"03AC",
      x"03B2", x"03B9", x"03C0", x"03C6", x"03CD", x"03D3", x"03DA", x"03E0", x"03E7", x"03ED", x"03F4", x"03FA", x"0401", x"0407", x"040E", x"0414",
      x"041B", x"0422", x"0428", x"042E", x"0435", x"043C", x"0442", x"0449", x"044F", x"0456", x"045C", x"0463", x"0469", x"0470", x"0476", x"047D",
      x"0484", x"048A", x"0490", x"0497", x"049E", x"04A4", x"04AB", x"04B1", x"04B8", x"04BE", x"04C5", x"04CB", x"04D2", x"04D8", x"04DF", x"04E5",
      x"04EC", x"04F2", x"04F9", x"0500", x"0506", x"050D", x"0513", x"051A", x"0520", x"0527", x"052D", x"0534", x"053A", x"0541", x"0547", x"054E",
      x"0554", x"055B", x"0562", x"0568", x"056E", x"0575", x"057C", x"0582", x"0589", x"058F", x"0596", x"059C", x"05A3", x"05A9", x"05B0", x"05B6",
      x"05BD", x"05C4", x"05CA", x"05D0", x"05D7", x"05DE", x"05E4", x"05EB", x"05F1", x"05F8", x"05FE", x"0605", x"060B", x"0612", x"0618", x"061F",
      x"0625", x"062C", x"0632", x"0639", x"0640", x"0646", x"064C", x"0653", x"065A", x"0660", x"0667", x"066D", x"0674", x"067A", x"0681", x"0687",
      x"068E", x"0694", x"069B", x"06A2", x"06A8", x"06AE", x"06B5", x"06BC", x"06C2", x"06C9", x"06CF", x"06D6", x"06DC", x"06E3", x"06E9", x"06F0",
      x"06F6", x"06FD", x"0703", x"070A", x"0710", x"0717", x"071E", x"0724", x"072B", x"0731", x"0738", x"073E", x"0745", x"074B", x"0752", x"0758",
      x"075F", x"0765", x"076C", x"0772", x"0779", x"0780", x"0786", x"078C", x"0793", x"079A", x"07A0", x"07A7", x"07AD", x"07B4", x"07BA", x"07C1",
      x"07C7", x"07CE", x"07D4", x"07DB", x"07E1", x"07E8", x"07EE", x"07F5", x"07FC", x"0802", x"0809", x"080F", x"0816", x"081C", x"0823", x"0829",
      x"0830", x"0836", x"083D", x"0843", x"084A", x"0850", x"0857", x"085E", x"0864", x"086A", x"0871", x"0878", x"087E", x"0885", x"088B", x"0892",
      x"0898", x"089F", x"08A5", x"08AC", x"08B2", x"08B9", x"08C0", x"08C6", x"08CC", x"08D3", x"08DA", x"08E0", x"08E7", x"08ED", x"08F4", x"08FA",
      x"0901", x"0907", x"090E", x"0914", x"091B", x"0921", x"0928", x"092E", x"0935", x"093C", x"0942", x"0948", x"094F", x"0956", x"095C", x"0963",
      x"0969", x"0970", x"0976", x"097D", x"0983", x"098A", x"0990", x"0997", x"099E", x"09A4", x"09AA", x"09B1", x"09B8", x"09BE", x"09C5", x"09CB",
      x"09D2", x"09D8", x"09DF", x"09E5", x"09EC", x"09F2", x"09F9", x"09FF", x"0A06", x"0A0C", x"0A13", x"0A1A", x"0A20", x"0A26", x"0A2D", x"0A34",
      x"0A3A", x"0A41", x"0A47", x"0A4E", x"0A54", x"0A5B", x"0A61", x"0A68", x"0A6E", x"0A75", x"0A7C", x"0A82", x"0A88", x"0A8F", x"0A96", x"0A9C",
      x"0AA3", x"0AA9", x"0AB0", x"0AB6", x"0ABD", x"0AC3", x"0ACA", x"0AD0", x"0AD7", x"0ADD", x"0AE4", x"0AEA", x"0AF1", x"0AF8", x"0AFE", x"0B04",
      x"0B0B", x"0B12", x"0B18", x"0B1F", x"0B25", x"0B2C", x"0B32", x"0B39", x"0B3F", x"0B46", x"0B4C", x"0B53", x"0B5A", x"0B60", x"0B66", x"0B6D",
      x"0B74", x"0B7A", x"0B81", x"0B87", x"0B8E", x"0B94", x"0B9B", x"0BA1", x"0BA8", x"0BAE", x"0BB5", x"0BBB", x"0BC2", x"0BC8", x"0BCF", x"0BD6",
      x"0BDC", x"0BE2", x"0BE9", x"0BF0", x"0BF6", x"0BFD", x"0C03", x"0C0A", x"0C10", x"0C17", x"0C1D", x"0C24", x"0C2A", x"0C31", x"0C38", x"0C3E",
      x"0C44", x"0C4B", x"0C52", x"0C58", x"0C5F", x"0C65", x"0C6C", x"0C72", x"0C79", x"0C7F", x"0C86", x"0C8C", x"0C93", x"0C99", x"0CA0", x"0CA6",
      x"0CAD", x"0CB4", x"0CBA", x"0CC0", x"0CC7", x"0CCE", x"0CD4", x"0CDB", x"0CE1", x"0CE8", x"0CEE", x"0CF5", x"0CFB", x"0D02", x"0D08", x"0D0F",
      x"0D15", x"0D1C", x"0D22", x"0D29", x"0D30", x"0D36", x"0D3D", x"0D43", x"0D4A", x"0D50", x"0D57", x"0D5D", x"0D64", x"0D6A", x"0D71", x"0D77",
      x"0D7E", x"0D84", x"0D8B", x"0D92", x"0D98", x"0D9E", x"0DA5", x"0DAC", x"0DB2", x"0DB9", x"0DBF", x"0DC6", x"0DCC", x"0DD3", x"0DD9", x"0DE0",
      x"0DE6", x"0DED", x"0DF3", x"0DFA", x"0E00", x"0E07", x"0E0E", x"0E14", x"0E1A", x"0E21", x"0E28", x"0E2E", x"0E35", x"0E3B", x"0E42", x"0E48",
      x"0E4F", x"0E55", x"0E5C", x"0E62", x"0E69", x"0E70", x"0E76", x"0E7C", x"0E83", x"0E8A", x"0E90", x"0E97", x"0E9D", x"0EA4", x"0EAA", x"0EB1",
      x"0EB7", x"0EBE", x"0EC4", x"0ECB", x"0ED1", x"0ED8", x"0EDE", x"0EE5", x"0EEC", x"0EF2", x"0EF8", x"0EFF", x"0F06", x"0F0C", x"0F13", x"0F19",
      x"0F20", x"0F26", x"0F2D", x"0F33", x"0F3A", x"0F40", x"0F47", x"0F4D", x"0F54", x"0F5A", x"0F61", x"0F68", x"0F6E", x"0F74", x"0F7B", x"0F82",
      x"0F88", x"0F8F", x"0F95", x"0F9C", x"0FA2", x"0FA9", x"0FAF", x"0FB6", x"0FBC", x"0FC3", x"0FCA", x"0FD0", x"0FD6", x"0FDD", x"0FE4", x"0FEA",
      x"0FF1", x"0FF7", x"0FFE", x"1004", x"100B", x"1011", x"1018", x"101E", x"1025", x"102B", x"1032", x"1038", x"103F", x"1046", x"104C", x"1052",
      x"1059", x"1060", x"1066", x"106D", x"1073", x"107A", x"1080", x"1087", x"108D", x"1094", x"109A", x"10A1", x"10A7", x"10AE", x"10B4", x"10BB",
      x"10C2", x"10C8", x"10CE", x"10D5", x"10DC", x"10E2", x"10E9", x"10EF", x"10F6", x"10FC", x"1103", x"1109", x"1110", x"1116", x"111D", x"1123",
      x"112A", x"1130", x"1137", x"113E", x"1144", x"114B", x"1151", x"1158", x"115E", x"1165", x"116B", x"1172", x"1178", x"117F", x"1185", x"118C",
      x"1192", x"1199", x"11A0", x"11A6", x"11AC", x"11B3", x"11BA", x"11C0", x"11C7", x"11CD", x"11D4", x"11DA", x"11E1", x"11E7", x"11EE", x"11F4",
      x"11FB", x"1201", x"1208", x"120E", x"1215", x"121C", x"1222", x"1228", x"122F", x"1236", x"123C", x"1243", x"1249", x"1250", x"1256", x"125D",
      x"1263", x"126A", x"1270", x"1277", x"127D", x"1284", x"128A", x"1291", x"1298", x"129E", x"12A4", x"12AB", x"12B2", x"12B8", x"12BF", x"12C5",
      x"12CC", x"12D2", x"12D9", x"12DF", x"12E6", x"12EC", x"12F3", x"12F9", x"1300", x"1306", x"130D", x"1314", x"131A", x"1320", x"1327", x"132E",
      x"1334", x"133B", x"1341", x"1348", x"134E", x"1355", x"135B", x"1362", x"1368", x"136F", x"1375", x"137C", x"1382", x"1389", x"1390", x"1396",
      x"139C", x"13A3", x"13AA", x"13B0", x"13B7", x"13BD", x"13C4", x"13CA", x"13D1", x"13D7", x"13DE", x"13E4", x"13EB", x"13F1", x"13F8", x"13FE",
      x"1405", x"140C", x"1412", x"1418", x"141F", x"1426", x"142C", x"1433", x"1439", x"1440", x"1446", x"144D", x"1453", x"145A", x"1460", x"1467",
      x"146D", x"1474", x"147A", x"1481", x"1488", x"148E", x"1494", x"149B", x"14A2", x"14A8", x"14AF", x"14B5", x"14BC", x"14C2", x"14C9", x"14CF",
      x"14D6", x"14DC", x"14E3", x"14E9", x"14F0", x"14F6", x"14FD", x"1504", x"150A", x"1510", x"1517", x"151E", x"1524", x"152B", x"1531", x"1538",
      x"153E", x"1545", x"154B", x"1552", x"1558", x"155F", x"1565", x"156C", x"1572", x"1579", x"1580", x"1586", x"158C", x"1593", x"159A", x"15A0",
      x"15A7", x"15AD", x"15B4", x"15BA", x"15C1", x"15C7", x"15CE", x"15D4", x"15DB", x"15E1", x"15E8", x"15EE", x"15F5", x"15FC", x"1602", x"1608",
      x"160F", x"1616", x"161C", x"1623", x"1629", x"1630", x"1636", x"163D", x"1643", x"164A", x"1650", x"1657", x"165D", x"1664", x"166A", x"1671",
      x"1678", x"167E", x"1684", x"168B", x"1692", x"1698", x"169F", x"16A5", x"16AC", x"16B2", x"16B9", x"16BF", x"16C6", x"16CC", x"16D3", x"16D9",
      x"16E0", x"16E6", x"16ED", x"16F4", x"16FA", x"1700", x"1707", x"170E", x"1714", x"171B", x"1721", x"1728", x"172E", x"1735", x"173B", x"1742",
      x"1748", x"174F", x"1755", x"175C", x"1762", x"1769", x"1770", x"1776", x"177C", x"1783", x"178A", x"1790", x"1797", x"179D", x"17A4", x"17AA",
      x"17B1", x"17B7", x"17BE", x"17C4", x"17CB", x"17D1", x"17D8", x"17DE", x"17E5", x"17EC", x"17F2", x"17F8", x"17FF", x"1806", x"180C", x"1813",
      x"1819", x"1820", x"1826", x"182D", x"1833", x"183A", x"1840", x"1847", x"184D", x"1854", x"185A", x"1861", x"1867", x"186E", x"1874", x"187B",
      x"1882", x"1888", x"188E", x"1895", x"189C", x"18A2", x"18A9", x"18AF", x"18B6", x"18BC", x"18C3", x"18C9", x"18D0", x"18D6", x"18DD", x"18E3",
      x"18EA", x"18F0", x"18F7", x"18FE", x"1904", x"190A", x"1911", x"1918", x"191E", x"1925", x"192B", x"1932", x"1938", x"193F", x"1945", x"194C",
      x"1952", x"1959", x"195F", x"1966", x"196C", x"1973", x"197A", x"1980", x"1986", x"198D", x"1994", x"199A", x"19A1", x"19A7", x"19AE", x"19B4",
      x"19BB", x"19C1", x"19C8", x"19CE", x"19D5", x"19DB", x"19E2", x"19E8", x"19EF", x"19F5", x"19FC", x"1A02", x"1A09", x"1A10", x"1A16", x"1A1C",

      -- Config 3
      x"006E", x"006E", x"006E", x"006F", x"006F", x"006F", x"006F", x"006F", x"006F", x"006F", x"006F", x"006F", x"006F", x"006F", x"006F", x"006F",
      x"006F", x"006F", x"006F", x"006F", x"006F", x"006F", x"006F", x"006F", x"006F", x"006F", x"006F", x"0070", x"0070", x"0070", x"0070", x"0070",
      x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070",
      x"0070", x"0070", x"0070", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071",
      x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0072", x"0072", x"0072", x"0072", x"0072",
      x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072",
      x"0072", x"0072", x"0072", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073",
      x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0074", x"0074", x"0074", x"0074", x"0074",
      x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074",
      x"0074", x"0074", x"0074", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075",
      x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0076", x"0076", x"0076", x"0076", x"0076",
      x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076",
      x"0076", x"0076", x"0076", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077",
      x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0078", x"0078", x"0078", x"0078", x"0078",
      x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078",
      x"0078", x"0078", x"0078", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079",
      x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079",
      x"0079", x"007A", x"007A", x"007A", x"007A", x"007A", x"007A", x"007A", x"007A", x"007A", x"007B", x"007B", x"007B", x"007B", x"007B", x"007C",
      x"007C", x"007C", x"007C", x"007D", x"007D", x"007D", x"007D", x"007E", x"007E", x"007E", x"007F", x"007F", x"007F", x"0080", x"0080", x"0081",
      x"0081", x"0082", x"0082", x"0083", x"0083", x"0084", x"0084", x"0085", x"0085", x"0086", x"0086", x"0087", x"0088", x"0088", x"0089", x"008A",
      x"008A", x"008B", x"008C", x"008D", x"008D", x"008E", x"008F", x"0090", x"0091", x"0092", x"0093", x"0094", x"0095", x"0096", x"0097", x"0098",
      x"0099", x"009A", x"009B", x"009C", x"009D", x"009E", x"00A0", x"00A1", x"00A2", x"00A3", x"00A5", x"00A6", x"00A7", x"00A9", x"00AA", x"00AC",
      x"00AD", x"00AF", x"00B0", x"00B2", x"00B3", x"00B5", x"00B7", x"00B8", x"00BA", x"00BC", x"00BD", x"00BF", x"00C1", x"00C3", x"00C5", x"00C7",
      x"00C9", x"00CB", x"00CD", x"00CF", x"00D1", x"00D3", x"00D5", x"00D7", x"00D9", x"00DC", x"00DE", x"00E0", x"00E3", x"00E5", x"00E7", x"00EA",
      x"00EC", x"00EF", x"00F1", x"00F4", x"00F7", x"00F9", x"00FC", x"00FF", x"0101", x"0104", x"0107", x"010A", x"010D", x"0110", x"0113", x"0116",
      x"0119", x"011C", x"011F", x"0122", x"0126", x"0129", x"012C", x"0130", x"0133", x"0136", x"013A", x"013D", x"0141", x"0145", x"0148", x"014C",
      x"0150", x"0153", x"0157", x"015B", x"015F", x"0163", x"0167", x"016B", x"016F", x"0173", x"0177", x"017C", x"0180", x"0184", x"0189", x"018D",
      x"0191", x"0196", x"019A", x"019F", x"01A4", x"01A8", x"01AD", x"01B2", x"01B7", x"01BC", x"01C1", x"01C6", x"01CB", x"01D0", x"01D5", x"01DA",
      x"01DF", x"01E4", x"01EA", x"01EF", x"01F5", x"01FA", x"0200", x"0205", x"020B", x"0210", x"0216", x"021C", x"0222", x"0228", x"022E", x"0234",
      x"023A", x"0240", x"0246", x"024C", x"0252", x"0259", x"025F", x"0266", x"026C", x"0273", x"0279", x"0280", x"0287", x"028D", x"0294", x"029B",
      x"02A2", x"02A9", x"02B0", x"02B7", x"02BE", x"02C6", x"02CD", x"02D4", x"02DC", x"02E3", x"02EB", x"02F2", x"02FA", x"0302", x"0309", x"0311",
      x"0319", x"0321", x"0329", x"0331", x"0339", x"0342", x"034A", x"0352", x"035B", x"0363", x"036C", x"0374", x"037D", x"0385", x"038E", x"0397",
      x"021F", x"0222", x"0227", x"022C", x"0232", x"0238", x"023F", x"0246", x"024E", x"0255", x"025D", x"0266", x"026E", x"0277", x"0280", x"0289",
      x"0292", x"029B", x"02A5", x"02AF", x"02B9", x"02C3", x"02CD", x"02D7", x"02E2", x"02EC", x"02F7", x"0302", x"030D", x"0318", x"0323", x"032F",
      x"033A", x"0346", x"0351", x"035D", x"0369", x"0375", x"0381", x"038D", x"0399", x"03A6", x"03B2", x"03BF", x"03CB", x"03D8", x"03E5", x"03F2",
      x"03FF", x"040C", x"0419", x"0426", x"0433", x"0441", x"044E", x"045B", x"0469", x"0477", x"0484", x"0492", x"04A0", x"04AE", x"04BC", x"04CA",
      x"04D8", x"04E6", x"04F5", x"0503", x"0511", x"0520", x"052E", x"053D", x"054C", x"055A", x"0569", x"0578", x"0587", x"0596", x"05A5", x"05B4",
      x"05C3", x"05D2", x"05E1", x"05F0", x"0600", x"060F", x"061F", x"062E", x"063E", x"064D", x"065D", x"066D", x"067C", x"068C", x"069C", x"06AC",
      x"06BC", x"06CC", x"06DC", x"06EC", x"06FC", x"070D", x"071D", x"072D", x"073D", x"074E", x"075E", x"076F", x"077F", x"0790", x"07A1", x"07B1",
      x"07C2", x"07D3", x"07E4", x"07F4", x"0805", x"0816", x"0827", x"0838", x"0849", x"085B", x"086C", x"087D", x"088E", x"089F", x"08B1", x"08C2",
      x"08D4", x"08E5", x"08F7", x"0908", x"091A", x"092B", x"093D", x"094F", x"0960", x"0972", x"0984", x"0996", x"09A8", x"09BA", x"09CC", x"09DE",
      x"09F0", x"0A02", x"0A14", x"0A26", x"0A38", x"0A4A", x"0A5D", x"0A6F", x"0A81", x"0A94", x"0AA6", x"0AB8", x"0ACB", x"0ADD", x"0AF0", x"0B03",
      x"0B15", x"0B28", x"0B3B", x"0B4D", x"0B60", x"0B73", x"0B86", x"0B99", x"0BAB", x"0BBE", x"0BD1", x"0BE4", x"0BF7", x"0C0A", x"0C1D", x"0C31",
      x"0C44", x"0C57", x"0C6A", x"0C7D", x"0C91", x"0CA4", x"0CB7", x"0CCB", x"0CDE", x"0CF2", x"0D05", x"0D19", x"0D2C", x"0D40", x"0D53", x"0D67",
      x"0D7B", x"0D8E", x"0DA2", x"0DB6", x"0DCA", x"0DDE", x"0DF1", x"0E05", x"0E19", x"0E2D", x"0E41", x"0E55", x"0E69", x"0E7D", x"0E91", x"0EA5",
      x"0EBA", x"0ECE", x"0EE2", x"0EF6", x"0F0A", x"0F1F", x"0F33", x"0F47", x"0F5C", x"0F70", x"0F85", x"0F99", x"0FAE", x"0FC2", x"0FD7", x"0FEB",
      x"1000", x"1014", x"1029", x"103E", x"1052", x"106A", x"1080", x"1095", x"10AA", x"10BF", x"10D3", x"10E8", x"10FC", x"1110", x"1124", x"1138",
      x"114B", x"115F", x"1173", x"1186", x"1199", x"11AD", x"11C0", x"11D4", x"11E7", x"11FA", x"120D", x"1220", x"1233", x"1246", x"1259", x"126C",
      x"127F", x"1292", x"12A5", x"12B8", x"12CA", x"12DD", x"12F0", x"1302", x"1315", x"1328", x"133A", x"134D", x"135F", x"1372", x"1385", x"1397",
      x"13A9", x"13BC", x"13CE", x"13E1", x"13F3", x"1406", x"1418", x"142A", x"143D", x"144F", x"1461", x"1473", x"1486", x"1498", x"14AA", x"14BC",
      x"14CE", x"14E1", x"14F3", x"1505", x"1517", x"1529", x"153B", x"154D", x"155F", x"1571", x"1583", x"1595", x"15A7", x"15B9", x"15CB", x"15DD",
      x"15EF", x"1601", x"1613", x"1625", x"1637", x"1649", x"165B", x"166D", x"167F", x"1691", x"16A2", x"16B4", x"16C6", x"16D8", x"16EA", x"16FC",
      x"170D", x"171F", x"1731", x"1743", x"1754", x"1766", x"1778", x"178A", x"179B", x"17AD", x"17BF", x"17D0", x"17E2", x"17F4", x"1805", x"1817",
      x"1829", x"183A", x"184C", x"185E", x"186F", x"1881", x"1892", x"18A4", x"18B6", x"18C7", x"18D9", x"18EA", x"18FC", x"190D", x"191F", x"1930",
      x"1942", x"1954", x"1965", x"1977", x"1988", x"199A", x"19AB", x"19BC", x"19CE", x"19DF", x"19F1", x"1A02", x"1A14", x"1A25", x"1A37", x"1A48",
      x"1A59", x"1A6B", x"1A7C", x"1A8E", x"1A9F", x"1AB0", x"1AC2", x"1AD3", x"1AE5", x"1AF6", x"1B07", x"1B19", x"1B2A", x"1B3B", x"1B4D", x"1B5E",
      x"1B6F", x"1B81", x"1B92", x"1BA3", x"1BB4", x"1BC6", x"1BD7", x"1BE8", x"1BFA", x"1C0B", x"1C1C", x"1C2D", x"1C3F", x"1C50", x"1C61", x"1C72",
      x"1C84", x"1C95", x"1CA6", x"1CB7", x"1CC8", x"1CDA", x"1CEB", x"1CFC", x"1D0D", x"1D1E", x"1D30", x"1D41", x"1D52", x"1D63", x"1D74", x"1D85",
      x"1D97", x"1DA8", x"1DB9", x"1DCA", x"1DDB", x"1DEC", x"1DFD", x"1E0F", x"1E20", x"1E31", x"1E42", x"1E53", x"1E64", x"1E75", x"1E86", x"1E97",
      x"1EA8", x"1EBA", x"1ECB", x"1EDC", x"1EED", x"1EFE", x"1F0F", x"1F20", x"1F31", x"1F42", x"1F53", x"1F64", x"1F75", x"1F86", x"1F97", x"1FA8",
      x"1FB9", x"1FCA", x"1FDB", x"1FEC", x"1FFD", x"200E", x"201F", x"2030", x"2041", x"2052", x"2063", x"2074", x"2085", x"2096", x"20A7", x"20B8",
      x"20C9", x"20DA", x"20EB", x"20FC", x"210D", x"211E", x"212F", x"213F", x"2150", x"2161", x"2172", x"2183", x"2194", x"21A5", x"21B6", x"21C7",
      x"21D8", x"21E9", x"21F9", x"220A", x"221B", x"222C", x"223D", x"224E", x"225F", x"2270", x"2280", x"2291", x"22A2", x"22B3", x"22C4", x"22D5",
      x"22E5", x"22F6", x"2307", x"2318", x"2329", x"233A", x"234A", x"235B", x"236C", x"237D", x"238E", x"239E", x"23AF", x"23C0", x"23D1", x"23E2",

      -- Config 4
      x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045",
      x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045",
      x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046",
      x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047",
      x"0047", x"0047", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0049", x"0049", x"0049", x"0049",
      x"0049", x"0049", x"0049", x"0049", x"004A", x"004A", x"004A", x"004A", x"004A", x"004A", x"004A", x"004A", x"004B", x"004B", x"004B", x"004B",
      x"004B", x"004B", x"004B", x"004C", x"004C", x"004C", x"004C", x"004C", x"004C", x"004C", x"004D", x"004D", x"004D", x"004D", x"004D", x"004D",
      x"004E", x"004E", x"004E", x"004E", x"004E", x"004E", x"004F", x"004F", x"004F", x"004F", x"004F", x"0050", x"0050", x"0050", x"0050", x"0050",
      x"0051", x"0051", x"0051", x"0051", x"0051", x"0052", x"0052", x"0052", x"0052", x"0052", x"0053", x"0053", x"0053", x"0053", x"0053", x"0054",
      x"0054", x"0054", x"0054", x"0055", x"0055", x"0055", x"0055", x"0055", x"0056", x"0056", x"0056", x"0056", x"0057", x"0057", x"0057", x"0057",
      x"0058", x"0058", x"0058", x"0058", x"0059", x"0059", x"0059", x"0059", x"005A", x"005A", x"005A", x"005A", x"005B", x"005B", x"005B", x"005C",
      x"005C", x"005C", x"005C", x"005D", x"005D", x"005D", x"005E", x"005E", x"005E", x"005E", x"005F", x"005F", x"005F", x"0060", x"0060", x"0060",
      x"0061", x"0061", x"0061", x"0061", x"0062", x"0062", x"0062", x"0063", x"0063", x"0063", x"0064", x"0064", x"0064", x"0065", x"0065", x"0065",
      x"0066", x"0066", x"0066", x"0067", x"0067", x"0067", x"0068", x"0068", x"0068", x"0069", x"0069", x"0069", x"006A", x"006A", x"006A", x"006B",
      x"006B", x"006C", x"006C", x"006C", x"006D", x"006D", x"006D", x"006E", x"006E", x"006F", x"006F", x"006F", x"0070", x"0070", x"0070", x"0071",
      x"0071", x"0072", x"0072", x"0072", x"0073", x"0073", x"0074", x"0074", x"0074", x"0075", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079",
      x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079",
      x"0079", x"007A", x"007A", x"007A", x"007A", x"007A", x"007A", x"007A", x"007A", x"007A", x"007B", x"007B", x"007B", x"007B", x"007B", x"007C",
      x"007C", x"007C", x"007C", x"007D", x"007D", x"007D", x"007D", x"007E", x"007E", x"007E", x"007F", x"007F", x"007F", x"0080", x"0080", x"0081",
      x"0081", x"0082", x"0082", x"0083", x"0083", x"0084", x"0084", x"0085", x"0085", x"0086", x"0086", x"0087", x"0088", x"0088", x"0089", x"008A",
      x"008A", x"008B", x"008C", x"008D", x"008D", x"008E", x"008F", x"0090", x"0091", x"0092", x"0093", x"0094", x"0095", x"0096", x"0097", x"0098",
      x"0099", x"009A", x"009B", x"009C", x"009D", x"009E", x"00A0", x"00A1", x"00A2", x"00A3", x"00A5", x"00A6", x"00A7", x"00A9", x"00AA", x"00AC",
      x"00AD", x"00AF", x"00B0", x"00B2", x"00B3", x"00B5", x"00B7", x"00B8", x"00BA", x"00BC", x"00BD", x"00BF", x"00C1", x"00C3", x"00C5", x"00C7",
      x"00C9", x"00CB", x"00CD", x"00CF", x"00D1", x"00D3", x"00D5", x"00D7", x"00D9", x"00DC", x"00DE", x"00E0", x"00E3", x"00E5", x"00E7", x"00EA",
      x"00EC", x"00EF", x"00F1", x"00F4", x"00F7", x"00F9", x"00FC", x"00FF", x"0101", x"0104", x"0107", x"010A", x"010D", x"0110", x"0113", x"0116",
      x"0119", x"011C", x"011F", x"0122", x"0126", x"0129", x"012C", x"0130", x"0133", x"0136", x"013A", x"013D", x"0141", x"0145", x"0148", x"014C",
      x"0150", x"0153", x"0157", x"015B", x"015F", x"0163", x"0167", x"016B", x"016F", x"0173", x"0177", x"017C", x"0180", x"0184", x"0189", x"018D",
      x"0191", x"0196", x"019A", x"019F", x"01A4", x"01A8", x"01AD", x"01B2", x"01B7", x"01BC", x"01C1", x"01C6", x"01CB", x"01D0", x"01D5", x"01DA",
      x"01DF", x"01E4", x"01EA", x"01EF", x"01F5", x"01FA", x"0200", x"0205", x"020B", x"0210", x"0216", x"021C", x"0222", x"0228", x"022E", x"0234",
      x"023A", x"0240", x"0246", x"024C", x"0252", x"0259", x"025F", x"0266", x"026C", x"0273", x"0279", x"0280", x"0287", x"028D", x"0294", x"029B",
      x"02A2", x"02A9", x"02B0", x"02B7", x"02BE", x"02C6", x"02CD", x"02D4", x"02DC", x"02E3", x"02EB", x"02F2", x"02FA", x"0302", x"0309", x"0311",
      x"0319", x"0321", x"0329", x"0331", x"0339", x"0342", x"034A", x"0352", x"035B", x"0363", x"036C", x"0374", x"037D", x"0385", x"038E", x"0397",
      x"021F", x"0222", x"0227", x"022C", x"0232", x"0238", x"023F", x"0246", x"024E", x"0255", x"025D", x"0266", x"026E", x"0277", x"0280", x"0289",
      x"0292", x"029B", x"02A5", x"02AF", x"02B9", x"02C3", x"02CD", x"02D7", x"02E2", x"02EC", x"02F7", x"0302", x"030D", x"0318", x"0323", x"032F",
      x"033A", x"0346", x"0351", x"035D", x"0369", x"0375", x"0381", x"038D", x"0399", x"03A6", x"03B2", x"03BF", x"03CB", x"03D8", x"03E5", x"03F2",
      x"03FF", x"040C", x"0419", x"0426", x"0433", x"0441", x"044E", x"045B", x"0469", x"0477", x"0484", x"0492", x"04A0", x"04AE", x"04BC", x"04CA",
      x"04D8", x"04E6", x"04F5", x"0503", x"0511", x"0520", x"052E", x"053D", x"054C", x"055A", x"0569", x"0578", x"0587", x"0596", x"05A5", x"05B4",
      x"05C3", x"05D2", x"05E1", x"05F0", x"0600", x"060F", x"061F", x"062E", x"063E", x"064D", x"065D", x"066D", x"067C", x"068C", x"069C", x"06AC",
      x"06BC", x"06CC", x"06DC", x"06EC", x"06FC", x"070D", x"071D", x"072D", x"073D", x"074E", x"075E", x"076F", x"077F", x"0790", x"07A1", x"07B1",
      x"07C2", x"07D3", x"07E4", x"07F4", x"0805", x"0816", x"0827", x"0838", x"0849", x"085B", x"086C", x"087D", x"088E", x"089F", x"08B1", x"08C2",
      x"08D4", x"08E5", x"08F7", x"0908", x"091A", x"092B", x"093D", x"094F", x"0960", x"0972", x"0984", x"0996", x"09A8", x"09BA", x"09CC", x"09DE",
      x"09F0", x"0A02", x"0A14", x"0A26", x"0A38", x"0A4A", x"0A5D", x"0A6F", x"0A81", x"0A94", x"0AA6", x"0AB8", x"0ACB", x"0ADD", x"0AF0", x"0B03",
      x"0B15", x"0B28", x"0B3B", x"0B4D", x"0B60", x"0B73", x"0B86", x"0B99", x"0BAB", x"0BBE", x"0BD1", x"0BE4", x"0BF7", x"0C0A", x"0C1D", x"0C31",
      x"0C44", x"0C57", x"0C6A", x"0C7D", x"0C91", x"0CA4", x"0CB7", x"0CCB", x"0CDE", x"0CF2", x"0D05", x"0D19", x"0D2C", x"0D40", x"0D53", x"0D67",
      x"0D7B", x"0D8E", x"0DA2", x"0DB6", x"0DCA", x"0DDE", x"0DF1", x"0E05", x"0E19", x"0E2D", x"0E41", x"0E55", x"0E69", x"0E7D", x"0E91", x"0EA5",
      x"0EBA", x"0ECE", x"0EE2", x"0EF6", x"0F0A", x"0F1F", x"0F33", x"0F47", x"0F5C", x"0F70", x"0F85", x"0F99", x"0FAE", x"0FC2", x"0FD7", x"0FEB",
      x"1000", x"1014", x"1029", x"103E", x"1052", x"1068", x"107A", x"108A", x"109A", x"10A8", x"10B7", x"10C5", x"10D3", x"10E0", x"10EE", x"10FB",
      x"1108", x"1114", x"1121", x"112D", x"113A", x"1146", x"1152", x"115E", x"116A", x"1176", x"1182", x"118D", x"1199", x"11A4", x"11B0", x"11BB",
      x"11C7", x"11D2", x"11DD", x"11E8", x"11F3", x"11FE", x"1209", x"1214", x"121F", x"122A", x"1235", x"1240", x"124A", x"1255", x"1260", x"126A",
      x"1275", x"127F", x"128A", x"1294", x"129F", x"12A9", x"12B4", x"12BE", x"12C8", x"12D3", x"12DD", x"12E7", x"12F1", x"12FB", x"1306", x"1310",
      x"131A", x"1324", x"132E", x"1338", x"1342", x"134C", x"1356", x"1360", x"136A", x"1373", x"137D", x"1387", x"1391", x"139B", x"13A5", x"13AE",
      x"13B8", x"13C2", x"13CB", x"13D5", x"13DF", x"13E8", x"13F2", x"13FC", x"1405", x"140F", x"1418", x"1422", x"142B", x"1435", x"143E", x"1448",
      x"1451", x"145B", x"1464", x"146E", x"1477", x"1480", x"148A", x"1493", x"149C", x"14A6", x"14AF", x"14B8", x"14C2", x"14CB", x"14D4", x"14DD",
      x"14E7", x"14F0", x"14F9", x"1502", x"150B", x"1515", x"151E", x"1527", x"1530", x"1539", x"1542", x"154B", x"1554", x"155E", x"1567", x"1570",
      x"1579", x"1582", x"158B", x"1594", x"159D", x"15A6", x"15AF", x"15B8", x"15C1", x"15CA", x"15D2", x"15DB", x"15E4", x"15ED", x"15F6", x"15FF",
      x"1608", x"1611", x"161A", x"1622", x"162B", x"1634", x"163D", x"1646", x"164F", x"1657", x"1660", x"1669", x"1672", x"167A", x"1683", x"168C",
      x"1695", x"169D", x"16A6", x"16AF", x"16B8", x"16C0", x"16C9", x"16D2", x"16DA", x"16E3", x"16EC", x"16F4", x"16FD", x"1705", x"170E", x"1717",
      x"171F", x"1728", x"1730", x"1739", x"1742", x"174A", x"1753", x"175B", x"1764", x"176C", x"1775", x"177D", x"1786", x"178E", x"1797", x"179F",
      x"17A8", x"17B0", x"17B9", x"17C1", x"17CA", x"17D2", x"17DB", x"17E3", x"17EC", x"17F4", x"17FC", x"1805", x"180D", x"1816", x"181E", x"1827",
      x"182F", x"1837", x"1840", x"1848", x"1850", x"1859", x"1861", x"1869", x"1872", x"187A", x"1882", x"188B", x"1893", x"189B", x"18A4", x"18AC",
      x"18B4", x"18BD", x"18C5", x"18CD", x"18D5", x"18DE", x"18E6", x"18EE", x"18F6", x"18FF", x"1907", x"190F", x"1917", x"1920", x"1928", x"1930",
      x"1938", x"1940", x"1949", x"1951", x"1959", x"1961", x"1969", x"1971", x"197A", x"1982", x"198A", x"1992", x"199A", x"19A2", x"19AA", x"19B3",
      x"19BB", x"19C3", x"19CB", x"19D3", x"19DB", x"19E3", x"19EB", x"19F3", x"19FC", x"1A04", x"1A0C", x"1A14", x"1A1C", x"1A24", x"1A2C", x"1A34",
      x"1A3C", x"1A44", x"1A4C", x"1A54", x"1A5C", x"1A64", x"1A6C", x"1A74", x"1A7C", x"1A84", x"1A8C", x"1A94", x"1A9C", x"1AA4", x"1AAC", x"1AB4",

      -- Config 5
      x"007A", x"007A", x"007A", x"007A", x"007A", x"007A", x"007B", x"007B", x"007B", x"007B", x"007B", x"007B", x"007B", x"007C", x"007C", x"007C",
      x"007C", x"007C", x"007C", x"007C", x"007C", x"007C", x"007C", x"007C", x"007C", x"007C", x"007C", x"007C", x"007C", x"007D", x"007D", x"007D",
      x"007D", x"007D", x"007D", x"007D", x"007E", x"007E", x"007E", x"007E", x"007E", x"007E", x"007E", x"007E", x"007E", x"007E", x"007E", x"007E",
      x"007E", x"007E", x"007E", x"007F", x"007F", x"007F", x"007F", x"007F", x"007F", x"007F", x"007F", x"0080", x"0080", x"0080", x"0080", x"0080",
      x"0080", x"0080", x"0080", x"0080", x"0080", x"0081", x"0081", x"0081", x"0081", x"0081", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082",
      x"0082", x"0083", x"0083", x"0083", x"0083", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0085", x"0085", x"0085", x"0085",
      x"0085", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0087", x"0087", x"0087", x"0087", x"0088", x"0088", x"0088", x"0088",
      x"0088", x"0088", x"0088", x"0089", x"0089", x"0089", x"0089", x"0089", x"008A", x"008A", x"008A", x"008A", x"008A", x"008A", x"008A", x"008B",
      x"008B", x"008C", x"008C", x"008C", x"008C", x"008D", x"008E", x"008E", x"008E", x"008F", x"008F", x"0090", x"0090", x"0090", x"0091", x"0092",
      x"0092", x"0092", x"0093", x"0093", x"0094", x"0094", x"0094", x"0095", x"0096", x"0096", x"0096", x"0097", x"0097", x"0098", x"0098", x"0098",
      x"0099", x"009A", x"009A", x"009A", x"009A", x"009B", x"009C", x"009C", x"009C", x"009D", x"009D", x"009E", x"009E", x"009E", x"009F", x"009F",
      x"00A0", x"00A0", x"00A1", x"00A1", x"00A2", x"00A2", x"00A2", x"00A3", x"00A3", x"00A4", x"00A4", x"00A5", x"00A5", x"00A6", x"00A6", x"00A6",
      x"00A7", x"00A8", x"00A9", x"00AA", x"00AB", x"00AC", x"00AD", x"00AE", x"00AF", x"00B0", x"00B1", x"00B2", x"00B4", x"00B4", x"00B6", x"00B6",
      x"00B8", x"00B8", x"00BA", x"00BA", x"00BC", x"00BD", x"00BE", x"00BF", x"00C0", x"00C1", x"00C2", x"00C3", x"00C4", x"00C5", x"00C6", x"00C7",
      x"00C8", x"00C9", x"00CA", x"00CC", x"00CC", x"00CE", x"00CE", x"00D0", x"00D0", x"00D2", x"00D2", x"00D4", x"00D5", x"00D6", x"00D7", x"00D8",
      x"00D9", x"00DA", x"00DB", x"00DC", x"00DD", x"00DE", x"00DF", x"00E0", x"00E1", x"00E2", x"00E4", x"00E4", x"00E6", x"00E6", x"00E8", x"00E8",
      x"00EA", x"00ED", x"00F0", x"00F3", x"00F6", x"00FA", x"00FC", x"0100", x"0103", x"0106", x"0109", x"010C", x"010F", x"0112", x"0116", x"0119",
      x"011C", x"011F", x"0122", x"0125", x"0128", x"012C", x"012E", x"0132", x"0135", x"0138", x"013B", x"013E", x"0142", x"0144", x"0148", x"014B",
      x"014E", x"0151", x"0154", x"0158", x"015A", x"015E", x"0161", x"0164", x"0167", x"016A", x"016E", x"0170", x"0174", x"0177", x"017A", x"017D",
      x"0180", x"0183", x"0186", x"018A", x"018D", x"0190", x"0193", x"0196", x"0199", x"019C", x"01A0", x"01A3", x"01A6", x"01A9", x"01AC", x"01AF",
      x"01B2", x"01BA", x"01C1", x"01C8", x"01CF", x"01D6", x"01DD", x"01E4", x"01EC", x"01F2", x"01FA", x"0201", x"0208", x"020F", x"0216", x"021E",
      x"0225", x"022C", x"0233", x"023A", x"0241", x"0248", x"0250", x"0256", x"025E", x"0265", x"026C", x"0273", x"027A", x"0282", x"0289", x"0290",
      x"0297", x"029E", x"02A5", x"02AC", x"02B4", x"02BA", x"02C2", x"02C9", x"02D0", x"02D7", x"02DE", x"02E6", x"02ED", x"02F4", x"02FB", x"0302",
      x"0309", x"0310", x"0318", x"031E", x"0326", x"032D", x"0334", x"033B", x"0342", x"034A", x"0351", x"0358", x"035F", x"0366", x"036E", x"0374",
      x"037C", x"0388", x"0394", x"03A0", x"03AC", x"03B8", x"03C5", x"03D1", x"03DD", x"03EA", x"03F6", x"0402", x"040E", x"041A", x"0426", x"0433",
      x"043F", x"044B", x"0457", x"0464", x"0470", x"047C", x"0488", x"0494", x"04A0", x"04AD", x"04B9", x"04C5", x"04D2", x"04DE", x"04EA", x"04F6",
      x"0502", x"0512", x"0522", x"0532", x"0541", x"0551", x"0560", x"0570", x"0580", x"0590", x"059F", x"05AF", x"05BF", x"05CE", x"05DE", x"05EE",
      x"05FE", x"060E", x"061D", x"062D", x"063C", x"064C", x"065C", x"066C", x"067C", x"068B", x"069B", x"06AA", x"06BA", x"06CA", x"06DA", x"06EA",
      x"06F9", x"070C", x"0720", x"0733", x"0746", x"075A", x"076D", x"0780", x"0793", x"07A6", x"07BA", x"07CD", x"07E0", x"07F4", x"0806", x"081A",
      x"082D", x"0840", x"0854", x"0867", x"087A", x"088E", x"08A1", x"08B4", x"08C7", x"08DA", x"08EE", x"0901", x"0914", x"0928", x"093B", x"094E",
      x"0962", x"097A", x"0993", x"09AB", x"09C4", x"09DC", x"09F5", x"0A0E", x"0A26", x"0A3F", x"0A57", x"0A70", x"0A88", x"0AA1", x"0ABA", x"0AD2",
      x"0AEB", x"0B07", x"0B23", x"0B3F", x"0B5C", x"0B78", x"0B94", x"0BB0", x"0BCC", x"0BF6", x"0C20", x"0C4B", x"0C75", x"0CA6", x"0CD6", x"0D06",
      x"0A0A", x"0A26", x"0A42", x"0A5E", x"0A7A", x"0A92", x"0AA9", x"0AC1", x"0AD8", x"0AF0", x"0B07", x"0B1E", x"0B36", x"0B4D", x"0B65", x"0B7C",
      x"0B94", x"0BAC", x"0BC5", x"0BDE", x"0BF6", x"0C0F", x"0C28", x"0C40", x"0C59", x"0C72", x"0C8A", x"0CA3", x"0CBC", x"0CD4", x"0CED", x"0D06",
      x"0D1E", x"0D34", x"0D49", x"0D5E", x"0D73", x"0D88", x"0D9E", x"0DB3", x"0DC8", x"0DDD", x"0DF2", x"0E08", x"0E1D", x"0E32", x"0E47", x"0E5C",
      x"0E72", x"0E87", x"0E9C", x"0EB2", x"0EC7", x"0EDC", x"0EF1", x"0F06", x"0F1C", x"0F31", x"0F46", x"0F5C", x"0F71", x"0F86", x"0F9C", x"0FB1",
      x"0FC6", x"0FDB", x"0FEF", x"1004", x"1018", x"102C", x"1041", x"1055", x"106A", x"107E", x"1092", x"10A7", x"10BC", x"10D0", x"10E4", x"10F9",
      x"110E", x"1122", x"1136", x"114B", x"1160", x"1174", x"1188", x"119D", x"11B2", x"11C6", x"11DA", x"11EF", x"1204", x"1218", x"122D", x"1241",
      x"1256", x"126A", x"127F", x"1294", x"12A8", x"12BD", x"12D1", x"12E6", x"12FA", x"130F", x"1324", x"1338", x"134D", x"1362", x"1376", x"138B",
      x"13A0", x"13B4", x"13C9", x"13DE", x"13F2", x"1406", x"141B", x"1430", x"1445", x"145A", x"146E", x"1483", x"1498", x"14AC", x"14C1", x"14D6",
      x"14EA", x"1501", x"1518", x"152E", x"1544", x"155B", x"1572", x"1588", x"159F", x"15B6", x"15CC", x"15E2", x"15F9", x"1610", x"1626", x"163D",
      x"1654", x"166A", x"1681", x"1698", x"16AE", x"16C5", x"16DC", x"16F2", x"1709", x"1720", x"1736", x"174D", x"1764", x"177A", x"1791", x"17A8",
      x"17BF", x"17D6", x"17EC", x"1803", x"181A", x"1831", x"1848", x"185E", x"1875", x"188C", x"18A3", x"18BA", x"18D0", x"18E8", x"18FE", x"1915",
      x"192C", x"1943", x"195A", x"1970", x"1988", x"199E", x"19B6", x"19CC", x"19E3", x"19FA", x"1A11", x"1A28", x"1A3F", x"1A56", x"1A6D", x"1A84",
      x"1A9B", x"1AB2", x"1AC9", x"1AE0", x"1AF8", x"1B0E", x"1B26", x"1B3C", x"1B54", x"1B6B", x"1B82", x"1B99", x"1BB0", x"1BC7", x"1BDE", x"1BF6",
      x"1C0C", x"1C24", x"1C3B", x"1C52", x"1C6A", x"1C80", x"1C98", x"1CAF", x"1CC6", x"1CDE", x"1CF5", x"1D0C", x"1D24", x"1D3A", x"1D52", x"1D6A",
      x"1D80", x"1D98", x"1DAF", x"1DC7", x"1DDE", x"1DF6", x"1E0D", x"1E24", x"1E3C", x"1E53", x"1E6A", x"1E82", x"1E9A", x"1EB1", x"1EC8", x"1EE0",
      x"1EF7", x"1F0F", x"1F26", x"1F3E", x"1F55", x"1F6D", x"1F84", x"1F9C", x"1FB4", x"1FCB", x"1FE3", x"1FFA", x"2012", x"202A", x"2041", x"2059",
      x"2070", x"207F", x"208D", x"209B", x"20AA", x"20B8", x"20C6", x"20D4", x"20E2", x"20F0", x"20FF", x"210D", x"211C", x"212A", x"2138", x"2146",
      x"2154", x"2163", x"2171", x"217F", x"218E", x"219C", x"21AA", x"21B8", x"21C7", x"21D5", x"21E4", x"21F2", x"2200", x"220E", x"221D", x"222B",
      x"223A", x"2248", x"2256", x"2264", x"2273", x"2281", x"2290", x"229E", x"22AC", x"22BB", x"22C9", x"22D8", x"22E6", x"22F4", x"2302", x"2311",
      x"2320", x"232E", x"233C", x"234B", x"2359", x"2368", x"2376", x"2384", x"2393", x"23A2", x"23B0", x"23BE", x"23CD", x"23DC", x"23EA", x"23F8",
      x"2407", x"2412", x"241C", x"2427", x"2432", x"243C", x"2447", x"2452", x"245C", x"2466", x"2472", x"247C", x"2487", x"2492", x"249C", x"24A7",
      x"24B2", x"24BC", x"24C7", x"24D2", x"24DC", x"24E7", x"24F2", x"24FC", x"2507", x"2512", x"251C", x"2527", x"2532", x"253C", x"2547", x"2552",
      x"255C", x"2567", x"2572", x"257D", x"2588", x"2592", x"259D", x"25A8", x"25B2", x"25BD", x"25C8", x"25D3", x"25DE", x"25E8", x"25F3", x"25FE",
      x"2608", x"2614", x"261E", x"2629", x"2634", x"263E", x"2649", x"2654", x"265F", x"266A", x"2674", x"267F", x"268A", x"2694", x"26A0", x"26AA",
      x"26B5", x"26BB", x"26C1", x"26C7", x"26CD", x"26D3", x"26D8", x"26DE", x"26E4", x"26EA", x"26F0", x"26F6", x"26FC", x"2702", x"2708", x"270E",
      x"2714", x"271A", x"2720", x"2726", x"272C", x"2731", x"2737", x"273D", x"2743", x"2749", x"274F", x"2755", x"275B", x"2760", x"2766", x"276C",
      x"2772", x"2778", x"277E", x"2784", x"278A", x"2790", x"2796", x"279C", x"27A2", x"27A8", x"27AE", x"27B4", x"27BA", x"27C0", x"27C6", x"27CC",
      x"27D2", x"27D8", x"27DD", x"27E3", x"27E9", x"27EF", x"27F5", x"27FB", x"2801", x"2807", x"280D", x"2813", x"2819", x"281F", x"2824", x"282B",
      x"2830", x"2834", x"2836", x"283A", x"283D", x"2840", x"2842", x"2846", x"2848", x"284C", x"284F", x"2852", x"2854", x"2858", x"285B", x"285E",
      x"2861", x"2864", x"2866", x"286A", x"286D", x"2870", x"2873", x"2876", x"2879", x"287C", x"287F", x"2882", x"2885", x"2888", x"288B", x"288E",
      x"2891", x"2894", x"2897", x"289A", x"289D", x"28A0", x"28A3", x"28A6", x"28A9", x"28AC", x"28AF", x"28B2", x"28B5", x"28B8", x"28BB", x"28BE",
      x"28C1", x"28C4", x"28C7", x"28CA", x"28CD", x"28D0", x"28D3", x"28D6", x"28D9", x"28DC", x"28DF", x"28E2", x"28E5", x"28E8", x"28EB", x"28EE",

      -- Config 6
      x"00B8", x"00B8", x"00B8", x"00B8", x"00B8", x"00B8", x"00B9", x"00B9", x"00B9", x"00B9", x"00B9", x"00B9", x"00B9", x"00BA", x"00BA", x"00BA",
      x"00BA", x"00BA", x"00BA", x"00BA", x"00BA", x"00BA", x"00BB", x"00BB", x"00BB", x"00BB", x"00BB", x"00BB", x"00BB", x"00BC", x"00BC", x"00BC",
      x"00BC", x"00BC", x"00BC", x"00BC", x"00BD", x"00BD", x"00BD", x"00BD", x"00BD", x"00BD", x"00BD", x"00BD", x"00BE", x"00BE", x"00BE", x"00BE",
      x"00BE", x"00BE", x"00BE", x"00BF", x"00BF", x"00BF", x"00BF", x"00BF", x"00BF", x"00BF", x"00BF", x"00C0", x"00C0", x"00C0", x"00C0", x"00C0",
      x"00C0", x"00C0", x"00C1", x"00C1", x"00C1", x"00C2", x"00C2", x"00C2", x"00C2", x"00C2", x"00C3", x"00C3", x"00C3", x"00C4", x"00C4", x"00C4",
      x"00C4", x"00C5", x"00C5", x"00C5", x"00C5", x"00C6", x"00C6", x"00C6", x"00C6", x"00C7", x"00C7", x"00C7", x"00C8", x"00C8", x"00C8", x"00C8",
      x"00C8", x"00C9", x"00C9", x"00C9", x"00CA", x"00CA", x"00CA", x"00CA", x"00CB", x"00CB", x"00CB", x"00CB", x"00CC", x"00CC", x"00CC", x"00CC",
      x"00CD", x"00CD", x"00CD", x"00CE", x"00CE", x"00CE", x"00CE", x"00CE", x"00CF", x"00CF", x"00CF", x"00D0", x"00D0", x"00D0", x"00D0", x"00D1",
      x"00D1", x"00D2", x"00D2", x"00D3", x"00D3", x"00D4", x"00D5", x"00D6", x"00D6", x"00D7", x"00D7", x"00D8", x"00D9", x"00D9", x"00DA", x"00DB",
      x"00DB", x"00DC", x"00DD", x"00DD", x"00DE", x"00DE", x"00DF", x"00E0", x"00E1", x"00E1", x"00E2", x"00E3", x"00E3", x"00E4", x"00E4", x"00E5",
      x"00E6", x"00E7", x"00E7", x"00E8", x"00E8", x"00E9", x"00EA", x"00EA", x"00EB", x"00EC", x"00EC", x"00ED", x"00EE", x"00EE", x"00EF", x"00EF",
      x"00F0", x"00F1", x"00F2", x"00F2", x"00F3", x"00F3", x"00F4", x"00F5", x"00F5", x"00F6", x"00F7", x"00F8", x"00F8", x"00F9", x"00F9", x"00FA",
      x"00FB", x"00FC", x"00FE", x"00FF", x"0101", x"0103", x"0104", x"0106", x"0107", x"0109", x"010A", x"010C", x"010E", x"010F", x"0111", x"0112",
      x"0114", x"0115", x"0117", x"0118", x"011A", x"011C", x"011D", x"011F", x"0120", x"0122", x"0123", x"0125", x"0127", x"0128", x"012A", x"012B",
      x"012D", x"012E", x"0130", x"0132", x"0133", x"0135", x"0136", x"0138", x"0139", x"013B", x"013C", x"013E", x"0140", x"0141", x"0143", x"0144",
      x"0146", x"0147", x"0149", x"014B", x"014C", x"014E", x"014F", x"0151", x"0152", x"0154", x"0156", x"0157", x"0159", x"015A", x"015C", x"015D",
      x"015F", x"0164", x"0169", x"016D", x"0172", x"0177", x"017B", x"0180", x"0185", x"0189", x"018E", x"0193", x"0197", x"019C", x"01A1", x"01A6",
      x"01AA", x"01AF", x"01B4", x"01B8", x"01BD", x"01C2", x"01C6", x"01CB", x"01D0", x"01D5", x"01D9", x"01DE", x"01E3", x"01E7", x"01EC", x"01F1",
      x"01F6", x"01FA", x"01FF", x"0204", x"0208", x"020D", x"0212", x"0216", x"021B", x"0220", x"0225", x"0229", x"022E", x"0233", x"0237", x"023C",
      x"0241", x"0245", x"024A", x"024F", x"0254", x"0258", x"025D", x"0262", x"0266", x"026B", x"0270", x"0275", x"0279", x"027E", x"0283", x"0287",
      x"028C", x"0297", x"02A2", x"02AC", x"02B7", x"02C2", x"02CC", x"02D7", x"02E2", x"02EC", x"02F7", x"0302", x"030D", x"0317", x"0322", x"032D",
      x"0338", x"0342", x"034D", x"0358", x"0362", x"036D", x"0378", x"0382", x"038D", x"0398", x"03A3", x"03AD", x"03B8", x"03C3", x"03CE", x"03D8",
      x"03E3", x"03EE", x"03F8", x"0403", x"040E", x"0418", x"0423", x"042E", x"0439", x"0443", x"044E", x"0459", x"0464", x"046E", x"0479", x"0484",
      x"048E", x"0499", x"04A4", x"04AE", x"04B9", x"04C4", x"04CF", x"04D9", x"04E4", x"04EF", x"04FA", x"0504", x"050F", x"051A", x"0525", x"052F",
      x"053A", x"054C", x"055E", x"0571", x"0583", x"0595", x"05A8", x"05BA", x"05CC", x"05DF", x"05F1", x"0603", x"0616", x"0628", x"063A", x"064D",
      x"065F", x"0671", x"0683", x"0696", x"06A8", x"06BA", x"06CD", x"06DF", x"06F1", x"0704", x"0716", x"0728", x"073B", x"074D", x"075F", x"0772",
      x"0784", x"079C", x"07B3", x"07CB", x"07E2", x"07FA", x"0811", x"0829", x"0841", x"0858", x"086F", x"0887", x"089F", x"08B6", x"08CE", x"08E5",
      x"08FD", x"0915", x"092C", x"0944", x"095B", x"0973", x"098A", x"09A2", x"09BA", x"09D1", x"09E9", x"0A00", x"0A18", x"0A30", x"0A47", x"0A5F",
      x"0A76", x"0A93", x"0AB0", x"0ACD", x"0AEA", x"0B07", x"0B24", x"0B40", x"0B5D", x"0B7A", x"0B97", x"0BB4", x"0BD1", x"0BEE", x"0C0A", x"0C27",
      x"0C44", x"0C61", x"0C7E", x"0C9B", x"0CB8", x"0CD5", x"0CF2", x"0D0F", x"0D2B", x"0D48", x"0D65", x"0D82", x"0D9F", x"0DBC", x"0DD9", x"0DF6",
      x"0E13", x"0E38", x"0E5D", x"0E81", x"0EA6", x"0ECB", x"0EF0", x"0F15", x"0F3A", x"0F5F", x"0F83", x"0FA8", x"0FCD", x"0FF2", x"1017", x"103C",
      x"1061", x"108B", x"10B5", x"10DF", x"110A", x"1134", x"115E", x"1188", x"11B2", x"11F2", x"1231", x"1271", x"12B0", x"12F9", x"1341", x"138A",
      x"0F0F", x"0F3A", x"0F64", x"0F8E", x"0FB8", x"0FDB", x"0FFE", x"1022", x"1045", x"1068", x"108B", x"10AE", x"10D1", x"10F4", x"1118", x"113B",
      x"115E", x"1183", x"11A8", x"11CD", x"11F2", x"1217", x"123C", x"1261", x"1286", x"12AB", x"12D0", x"12F5", x"131A", x"133F", x"1364", x"1389",
      x"13AE", x"13CE", x"13EE", x"140D", x"142D", x"144D", x"146D", x"148D", x"14AD", x"14CC", x"14EC", x"150C", x"152C", x"154C", x"156B", x"158B",
      x"15AB", x"15CB", x"15EB", x"160B", x"162B", x"164B", x"166A", x"168A", x"16AA", x"16CA", x"16EA", x"170A", x"172A", x"174A", x"176A", x"178A",
      x"17AA", x"17C9", x"17E7", x"1806", x"1824", x"1843", x"1862", x"1880", x"189F", x"18BE", x"18DC", x"18FB", x"191A", x"1939", x"1957", x"1976",
      x"1995", x"19B3", x"19D2", x"19F1", x"1A10", x"1A2E", x"1A4D", x"1A6C", x"1A8B", x"1AAA", x"1AC8", x"1AE7", x"1B06", x"1B25", x"1B44", x"1B62",
      x"1B81", x"1BA0", x"1BBF", x"1BDE", x"1BFD", x"1C1C", x"1C3A", x"1C59", x"1C78", x"1C97", x"1CB6", x"1CD5", x"1CF4", x"1D13", x"1D32", x"1D51",
      x"1D70", x"1D8F", x"1DAE", x"1DCD", x"1DEC", x"1E0A", x"1E29", x"1E49", x"1E68", x"1E87", x"1EA6", x"1EC5", x"1EE4", x"1F03", x"1F22", x"1F41",
      x"1F60", x"1F82", x"1FA4", x"1FC5", x"1FE7", x"2009", x"202B", x"204D", x"206F", x"2091", x"20B2", x"20D4", x"20F6", x"2118", x"213A", x"215C",
      x"217E", x"21A0", x"21C2", x"21E4", x"2206", x"2228", x"224A", x"226C", x"228E", x"22B0", x"22D2", x"22F4", x"2316", x"2338", x"235A", x"237D",
      x"239F", x"23C1", x"23E3", x"2405", x"2427", x"244A", x"246C", x"248E", x"24B0", x"24D2", x"24F5", x"2517", x"2539", x"255C", x"257E", x"25A0",
      x"25C2", x"25E5", x"2607", x"2629", x"264C", x"266E", x"2691", x"26B3", x"26D5", x"26F8", x"271A", x"273D", x"275F", x"2782", x"27A4", x"27C7",
      x"27E9", x"280C", x"282E", x"2851", x"2874", x"2896", x"28B9", x"28DB", x"28FE", x"2921", x"2943", x"2966", x"2988", x"29AB", x"29CE", x"29F1",
      x"2A13", x"2A36", x"2A59", x"2A7C", x"2A9F", x"2AC1", x"2AE4", x"2B07", x"2B2A", x"2B4D", x"2B70", x"2B93", x"2BB6", x"2BD8", x"2BFB", x"2C1F",
      x"2C41", x"2C64", x"2C87", x"2CAB", x"2CCE", x"2CF1", x"2D14", x"2D37", x"2D5A", x"2D7D", x"2DA0", x"2DC3", x"2DE7", x"2E0A", x"2E2D", x"2E50",
      x"2E73", x"2E97", x"2EBA", x"2EDD", x"2F00", x"2F24", x"2F47", x"2F6A", x"2F8E", x"2FB1", x"2FD5", x"2FF8", x"301B", x"303F", x"3062", x"3086",
      x"30A9", x"30BF", x"30D4", x"30E9", x"30FF", x"3114", x"3129", x"313F", x"3154", x"3169", x"317F", x"3194", x"31AA", x"31BF", x"31D4", x"31EA",
      x"31FF", x"3215", x"322A", x"323F", x"3255", x"326A", x"3280", x"3295", x"32AB", x"32C0", x"32D6", x"32EB", x"3300", x"3316", x"332C", x"3341",
      x"3357", x"336C", x"3382", x"3397", x"33AD", x"33C2", x"33D8", x"33ED", x"3403", x"3419", x"342E", x"3444", x"3459", x"346F", x"3484", x"349A",
      x"34B0", x"34C5", x"34DB", x"34F1", x"3506", x"351C", x"3532", x"3547", x"355D", x"3573", x"3588", x"359E", x"35B4", x"35CA", x"35DF", x"35F5",
      x"360B", x"361B", x"362B", x"363B", x"364B", x"365B", x"366B", x"367B", x"368B", x"369A", x"36AB", x"36BB", x"36CB", x"36DB", x"36EA", x"36FB",
      x"370B", x"371B", x"372B", x"373B", x"374B", x"375B", x"376B", x"377B", x"378B", x"379B", x"37AB", x"37BB", x"37CB", x"37DB", x"37EB", x"37FB",
      x"380B", x"381B", x"382C", x"383C", x"384C", x"385C", x"386C", x"387C", x"388C", x"389C", x"38AD", x"38BD", x"38CD", x"38DD", x"38ED", x"38FD",
      x"390D", x"391E", x"392E", x"393E", x"394E", x"395E", x"396E", x"397E", x"398F", x"399F", x"39AF", x"39BF", x"39CF", x"39DF", x"39F0", x"3A00",
      x"3A10", x"3A19", x"3A22", x"3A2B", x"3A34", x"3A3D", x"3A45", x"3A4E", x"3A57", x"3A60", x"3A69", x"3A72", x"3A7B", x"3A83", x"3A8C", x"3A95",
      x"3A9E", x"3AA7", x"3AB0", x"3AB9", x"3AC2", x"3ACA", x"3AD3", x"3ADC", x"3AE5", x"3AEE", x"3AF7", x"3B00", x"3B09", x"3B11", x"3B1A", x"3B23",
      x"3B2C", x"3B35", x"3B3E", x"3B47", x"3B50", x"3B59", x"3B61", x"3B6A", x"3B73", x"3B7C", x"3B85", x"3B8E", x"3B97", x"3BA0", x"3BA9", x"3BB2",
      x"3BBB", x"3BC4", x"3BCC", x"3BD5", x"3BDE", x"3BE7", x"3BF0", x"3BF9", x"3C02", x"3C0B", x"3C14", x"3C1D", x"3C26", x"3C2F", x"3C37", x"3C41",
      x"3C49", x"3C4E", x"3C52", x"3C57", x"3C5C", x"3C60", x"3C64", x"3C69", x"3C6D", x"3C72", x"3C77", x"3C7B", x"3C7F", x"3C84", x"3C89", x"3C8D",
      x"3C92", x"3C96", x"3C9A", x"3C9F", x"3CA4", x"3CA8", x"3CAD", x"3CB1", x"3CB6", x"3CBA", x"3CBF", x"3CC3", x"3CC8", x"3CCC", x"3CD1", x"3CD5",
      x"3CDA", x"3CDE", x"3CE3", x"3CE7", x"3CEC", x"3CF0", x"3CF5", x"3CF9", x"3CFE", x"3D02", x"3D07", x"3D0B", x"3D10", x"3D15", x"3D19", x"3D1D",
      x"3D22", x"3D27", x"3D2B", x"3D30", x"3D34", x"3D39", x"3D3D", x"3D42", x"3D46", x"3D4B", x"3D4F", x"3D54", x"3D58", x"3D5D", x"3D61", x"3D66",

      -- Config 7
      x"0114", x"0114", x"0114", x"0114", x"0114", x"0114", x"0115", x"0115", x"0115", x"0115", x"0115", x"0115", x"0115", x"0117", x"0117", x"0117",
      x"0117", x"0117", x"0117", x"0117", x"0117", x"0117", x"0118", x"0118", x"0118", x"0118", x"0118", x"0118", x"0118", x"011A", x"011A", x"011A",
      x"011A", x"011A", x"011A", x"011A", x"011B", x"011B", x"011B", x"011B", x"011B", x"011B", x"011B", x"011B", x"011D", x"011D", x"011D", x"011D",
      x"011D", x"011D", x"011D", x"011E", x"011E", x"011E", x"011E", x"011E", x"011E", x"011E", x"011E", x"0120", x"0120", x"0120", x"0120", x"0120",
      x"0120", x"0120", x"0121", x"0121", x"0121", x"0123", x"0123", x"0123", x"0123", x"0123", x"0124", x"0124", x"0124", x"0126", x"0126", x"0126",
      x"0126", x"0127", x"0127", x"0127", x"0127", x"0129", x"0129", x"0129", x"0129", x"012A", x"012A", x"012A", x"012C", x"012C", x"012C", x"012C",
      x"012C", x"012D", x"012D", x"012D", x"012F", x"012F", x"012F", x"012F", x"0130", x"0130", x"0130", x"0130", x"0132", x"0132", x"0132", x"0132",
      x"0133", x"0133", x"0133", x"0135", x"0135", x"0135", x"0135", x"0135", x"0136", x"0136", x"0136", x"0138", x"0138", x"0138", x"0138", x"0139",
      x"0139", x"013B", x"013B", x"013C", x"013C", x"013E", x"013F", x"0141", x"0141", x"0142", x"0142", x"0144", x"0145", x"0145", x"0147", x"0148",
      x"0148", x"014A", x"014B", x"014B", x"014D", x"014D", x"014E", x"0150", x"0151", x"0151", x"0153", x"0154", x"0154", x"0156", x"0156", x"0157",
      x"0159", x"015A", x"015A", x"015C", x"015C", x"015D", x"015F", x"015F", x"0160", x"0162", x"0162", x"0163", x"0165", x"0165", x"0166", x"0166",
      x"0168", x"0169", x"016B", x"016B", x"016C", x"016C", x"016E", x"016F", x"016F", x"0171", x"0172", x"0174", x"0174", x"0175", x"0175", x"0177",
      x"0178", x"017A", x"017D", x"017E", x"0181", x"0184", x"0186", x"0189", x"018A", x"018D", x"018F", x"0192", x"0195", x"0196", x"0199", x"019B",
      x"019E", x"019F", x"01A2", x"01A4", x"01A7", x"01AA", x"01AB", x"01AE", x"01B0", x"01B3", x"01B4", x"01B7", x"01BA", x"01BC", x"01BF", x"01C0",
      x"01C3", x"01C5", x"01C8", x"01CB", x"01CC", x"01CF", x"01D1", x"01D4", x"01D5", x"01D8", x"01DA", x"01DD", x"01E0", x"01E1", x"01E4", x"01E6",
      x"01E9", x"01EA", x"01ED", x"01F0", x"01F2", x"01F5", x"01F6", x"01F9", x"01FB", x"01FE", x"0201", x"0202", x"0205", x"0207", x"020A", x"020B",
      x"020E", x"0216", x"021D", x"0223", x"022B", x"0232", x"0238", x"0240", x"0247", x"024D", x"0255", x"025C", x"0262", x"026A", x"0271", x"0279",
      x"027F", x"0286", x"028E", x"0294", x"029B", x"02A3", x"02A9", x"02B0", x"02B8", x"02BF", x"02C5", x"02CD", x"02D4", x"02DA", x"02E2", x"02E9",
      x"02F1", x"02F7", x"02FE", x"0306", x"030C", x"0313", x"031B", x"0321", x"0328", x"0330", x"0337", x"033D", x"0345", x"034C", x"0352", x"035A",
      x"0361", x"0367", x"036F", x"0376", x"037E", x"0384", x"038B", x"0393", x"0399", x"03A0", x"03A8", x"03AF", x"03B5", x"03BD", x"03C4", x"03CA",
      x"03D2", x"03E2", x"03F3", x"0402", x"0412", x"0423", x"0432", x"0442", x"0453", x"0462", x"0472", x"0483", x"0493", x"04A2", x"04B3", x"04C3",
      x"04D4", x"04E3", x"04F3", x"0504", x"0513", x"0523", x"0534", x"0543", x"0553", x"0564", x"0574", x"0583", x"0594", x"05A4", x"05B5", x"05C4",
      x"05D4", x"05E5", x"05F4", x"0604", x"0615", x"0624", x"0634", x"0645", x"0655", x"0664", x"0675", x"0685", x"0696", x"06A5", x"06B5", x"06C6",
      x"06D5", x"06E5", x"06F6", x"0705", x"0715", x"0726", x"0736", x"0745", x"0756", x"0766", x"0777", x"0786", x"0796", x"07A7", x"07B7", x"07C6",
      x"07D7", x"07F2", x"080D", x"0829", x"0844", x"085F", x"087C", x"0897", x"08B2", x"08CE", x"08E9", x"0904", x"0921", x"093C", x"0957", x"0973",
      x"098E", x"09A9", x"09C4", x"09E1", x"09FC", x"0A17", x"0A33", x"0A4E", x"0A69", x"0A86", x"0AA1", x"0ABC", x"0AD8", x"0AF3", x"0B0E", x"0B2B",
      x"0B46", x"0B6A", x"0B8C", x"0BB0", x"0BD3", x"0BF7", x"0C19", x"0C3D", x"0C61", x"0C84", x"0CA6", x"0CCA", x"0CEE", x"0D11", x"0D35", x"0D57",
      x"0D7B", x"0D9F", x"0DC2", x"0DE6", x"0E08", x"0E2C", x"0E4F", x"0E73", x"0E97", x"0EB9", x"0EDD", x"0F00", x"0F24", x"0F48", x"0F6A", x"0F8E",
      x"0FB1", x"0FDC", x"1008", x"1033", x"105F", x"108A", x"10B6", x"10E0", x"110B", x"1137", x"1162", x"118E", x"11B9", x"11E5", x"120F", x"123A",
      x"1266", x"1291", x"12BD", x"12E8", x"1314", x"133F", x"136B", x"1396", x"13C0", x"13EC", x"1417", x"1443", x"146E", x"149A", x"14C5", x"14F1",
      x"151C", x"1554", x"158B", x"15C1", x"15F9", x"1630", x"1668", x"169F", x"16D7", x"170E", x"1744", x"177C", x"17B3", x"17EB", x"1822", x"185A",
      x"1891", x"18D0", x"190F", x"194E", x"198F", x"19CE", x"1A0D", x"1A4C", x"1A8B", x"1AEB", x"1B49", x"1BA9", x"1C08", x"1C75", x"1CE1", x"1D4F",
      x"1696", x"16D7", x"1716", x"1755", x"1794", x"17C8", x"17FD", x"1833", x"1867", x"189C", x"18D0", x"1905", x"1939", x"196E", x"19A4", x"19D8",
      x"1A0D", x"1A44", x"1A7C", x"1AB3", x"1AEB", x"1B22", x"1B5A", x"1B91", x"1BC9", x"1C00", x"1C38", x"1C6F", x"1CA7", x"1CDE", x"1D16", x"1D4D",
      x"1D85", x"1DB5", x"1DE5", x"1E13", x"1E43", x"1E73", x"1EA3", x"1ED3", x"1F03", x"1F32", x"1F62", x"1F92", x"1FC2", x"1FF2", x"2020", x"2050",
      x"2080", x"20B0", x"20E0", x"2110", x"2140", x"2170", x"219F", x"21CF", x"21FF", x"222F", x"225F", x"228F", x"22BF", x"22EF", x"231F", x"234F",
      x"237F", x"23AD", x"23DA", x"2409", x"2436", x"2464", x"2493", x"24C0", x"24EE", x"251D", x"254A", x"2578", x"25A7", x"25D5", x"2602", x"2631",
      x"265F", x"268C", x"26BB", x"26E9", x"2718", x"2745", x"2773", x"27A2", x"27D0", x"27FF", x"282C", x"285A", x"2889", x"28B7", x"28E6", x"2913",
      x"2941", x"2970", x"299E", x"29CD", x"29FB", x"2A2A", x"2A57", x"2A85", x"2AB4", x"2AE2", x"2B11", x"2B3F", x"2B6E", x"2B9C", x"2BCB", x"2BF9",
      x"2C28", x"2C56", x"2C85", x"2CB3", x"2CE2", x"2D0F", x"2D3D", x"2D6D", x"2D9C", x"2DCA", x"2DF9", x"2E27", x"2E56", x"2E84", x"2EB3", x"2EE1",
      x"2F10", x"2F43", x"2F76", x"2FA7", x"2FDA", x"300D", x"3040", x"3073", x"30A6", x"30D9", x"310B", x"313E", x"3171", x"31A4", x"31D7", x"320A",
      x"323D", x"3270", x"32A3", x"32D6", x"3309", x"333C", x"336F", x"33A2", x"33D5", x"3408", x"343B", x"346E", x"34A1", x"34D4", x"3507", x"353B",
      x"356E", x"35A1", x"35D4", x"3607", x"363A", x"366F", x"36A2", x"36D5", x"3708", x"373B", x"376F", x"37A2", x"37D5", x"380A", x"383D", x"3870",
      x"38A3", x"38D7", x"390A", x"393D", x"3972", x"39A5", x"39D9", x"3A0C", x"3A3F", x"3A74", x"3AA7", x"3ADB", x"3B0E", x"3B43", x"3B76", x"3BAA",
      x"3BDD", x"3C12", x"3C45", x"3C79", x"3CAE", x"3CE1", x"3D15", x"3D48", x"3D7D", x"3DB1", x"3DE4", x"3E19", x"3E4C", x"3E80", x"3EB5", x"3EE9",
      x"3F1C", x"3F51", x"3F85", x"3FBA", x"3FEE", x"4021", x"4056", x"408A", x"40BF", x"40F3", x"4128", x"415C", x"4191", x"41C4", x"41F8", x"422E",
      x"4261", x"4296", x"42CA", x"4300", x"4335", x"4369", x"439E", x"43D2", x"4407", x"443B", x"4470", x"44A4", x"44DA", x"450F", x"4543", x"4578",
      x"45AC", x"45E2", x"4617", x"464B", x"4680", x"46B6", x"46EA", x"471F", x"4755", x"4789", x"47BF", x"47F4", x"4828", x"485E", x"4893", x"48C9",
      x"48FD", x"491E", x"493E", x"495D", x"497E", x"499E", x"49BD", x"49DE", x"49FE", x"4A1D", x"4A3E", x"4A5E", x"4A7F", x"4A9E", x"4ABE", x"4ADF",
      x"4AFE", x"4B1F", x"4B3F", x"4B5E", x"4B7F", x"4B9F", x"4BC0", x"4BDF", x"4C00", x"4C20", x"4C41", x"4C60", x"4C80", x"4CA1", x"4CC2", x"4CE1",
      x"4D02", x"4D22", x"4D43", x"4D62", x"4D83", x"4DA3", x"4DC4", x"4DE3", x"4E04", x"4E25", x"4E45", x"4E66", x"4E85", x"4EA6", x"4EC6", x"4EE7",
      x"4F08", x"4F27", x"4F48", x"4F69", x"4F89", x"4FAA", x"4FCB", x"4FEA", x"500B", x"502C", x"504C", x"506D", x"508E", x"50AF", x"50CE", x"50EF",
      x"5110", x"5128", x"5140", x"5158", x"5170", x"5188", x"51A0", x"51B8", x"51D0", x"51E7", x"5200", x"5218", x"5230", x"5248", x"525F", x"5278",
      x"5290", x"52A8", x"52C0", x"52D8", x"52F0", x"5308", x"5320", x"5338", x"5350", x"5368", x"5380", x"5398", x"53B0", x"53C8", x"53E0", x"53F8",
      x"5410", x"5428", x"5442", x"545A", x"5472", x"548A", x"54A2", x"54BA", x"54D2", x"54EA", x"5503", x"551B", x"5533", x"554B", x"5563", x"557B",
      x"5593", x"55AD", x"55C5", x"55DD", x"55F5", x"560D", x"5625", x"563D", x"5656", x"566E", x"5686", x"569E", x"56B6", x"56CE", x"56E8", x"5700",
      x"5718", x"5725", x"5733", x"5740", x"574E", x"575B", x"5767", x"5775", x"5782", x"5790", x"579D", x"57AB", x"57B8", x"57C4", x"57D2", x"57DF",
      x"57ED", x"57FA", x"5808", x"5815", x"5823", x"582F", x"583C", x"584A", x"5857", x"5865", x"5872", x"5880", x"588D", x"5899", x"58A7", x"58B4",
      x"58C2", x"58CF", x"58DD", x"58EA", x"58F8", x"5905", x"5911", x"591F", x"592C", x"593A", x"5947", x"5955", x"5962", x"5970", x"597D", x"598B",
      x"5998", x"59A6", x"59B2", x"59BF", x"59CD", x"59DA", x"59E8", x"59F5", x"5A03", x"5A10", x"5A1E", x"5A2B", x"5A39", x"5A46", x"5A52", x"5A61",
      x"5A6D", x"5A75", x"5A7B", x"5A82", x"5A8A", x"5A90", x"5A96", x"5A9D", x"5AA3", x"5AAB", x"5AB2", x"5AB8", x"5ABE", x"5AC6", x"5ACD", x"5AD3",
      x"5ADB", x"5AE1", x"5AE7", x"5AEE", x"5AF6", x"5AFC", x"5B03", x"5B09", x"5B11", x"5B17", x"5B1E", x"5B24", x"5B2C", x"5B32", x"5B39", x"5B3F",
      x"5B47", x"5B4D", x"5B54", x"5B5A", x"5B62", x"5B68", x"5B6F", x"5B75", x"5B7D", x"5B83", x"5B8A", x"5B90", x"5B98", x"5B9F", x"5BA5", x"5BAB",
      x"5BB3", x"5BBA", x"5BC0", x"5BC8", x"5BCE", x"5BD5", x"5BDB", x"5BE3", x"5BE9", x"5BF0", x"5BF6", x"5BFE", x"5C04", x"5C0B", x"5C11", x"5C19"
    );

    signal filter_q     : signed(17 downto 0);
    signal filter_f     : signed(17 downto 0);
    signal input_sc     : signed(21 downto 0);
    signal xa           : signed(17 downto 0);
    signal xb           : signed(17 downto 0);
    signal sum_b        : signed(21 downto 0);
    signal sub_a        : signed(21 downto 0);
    signal sub_b        : signed(21 downto 0);
    signal x_reg        : signed(21 downto 0) := (others => '0');
    signal bp_reg       : signed(21 downto 0);
    signal hp_reg       : signed(21 downto 0);
    signal lp_reg       : signed(21 downto 0);
    signal temp_reg     : signed(21 downto 0);
    signal error        : std_logic := '0';
    signal program_cnt  : integer range 0 to 15;
    signal scale_cnt    : integer range 0 to 23;

    signal instruction  : std_logic_vector(7 downto 0);

    alias  xa_select    : std_logic is instruction(0);
    alias  xb_select    : std_logic is instruction(1);
    alias  sub_a_sel    : std_logic is instruction(2);
    alias  sub_b_sel    : std_logic is instruction(3);
    alias  sum_to_lp    : std_logic is instruction(4);
    alias  sum_to_bp    : std_logic is instruction(5);
    alias  sub_to_hp    : std_logic is instruction(6);
    alias  mult_enable  : std_logic is instruction(7);

    -- operations to execute the filter:
    -- lp        = (f * bp_reg) + lp_reg
    -- hp_reg    = input - lp - (q * bp_reg)
    -- bp        = (f * hp_reg) + bp_reg   
    -- bp_reg    = bp              
    -- lp_reg    = lp              

    -- x_reg     = f * bp_reg           -- 10000000 -- 80
    -- lp_reg    = x_reg + lp_reg       -- 00010010 -- 12
    -- q_contrib = q * bp_reg           -- 10000001 -- 81
    -- temp      = input - lp           -- 00000000 -- 00 (can be merged with previous!)
    -- hp_reg    = temp - q_contrib     -- 01001100 -- 4C
    -- x_reg     = f * hp_reg           -- 10000010 -- 82
    -- bp_reg    = x_reg + bp_reg       -- 00100000 -- 20

    type t_byte_array is array(natural range <>) of std_logic_vector(7 downto 0);
    constant c_program  : t_byte_array := (X"80", X"12", X"81", X"4C", X"82", X"20", X"00");

begin
    process(ld_clk)
    begin
        if rising_edge(ld_clk) then
            if(ld_wr = '1') then
                coef(5120+to_integer(unsigned(ld_addr))) <= signed(ld_data);
            end if;
        end if;
    end process;

    -- Derive the actual 'f' and 'q' parameters
    i_q_table: entity work.Q_table
    port map (
        Q_reg       => filt_res,
        filter_q    => filter_q ); -- 2.16 format

    process(clock)
    begin
        if rising_edge(clock) then
            if(enable = '1') then
                filter_f <= "00" & coef(to_integer(cfg & filt_co(10 downto 1)));
            else
                filter_f <= "001111111111111111";
            end if;
        end if;
    end process;

    input_sc <= shift_right(input, 1) & "0000";

    -- now perform the arithmetic
    xa    <= filter_f when xa_select='0' else filter_q;
    xb    <= bp_reg(21 downto 4) when xb_select='0' else hp_reg (21 downto 4);
    sum_b <= bp_reg   when xb_select='0' else lp_reg;
    sub_a <= input_sc when sub_a_sel='0' else temp_reg;
    sub_b <= lp_reg   when sub_b_sel='0' else x_reg;
    
    process(clock)
        variable x_result   : signed(35 downto 0);
        variable sum_result : signed(21 downto 0);
        variable sub_result : signed(21 downto 0);
    begin
        if rising_edge(clock) then
            x_result := xa * xb;
            if mult_enable='1' then
                x_reg <= x_result(33 downto 12);
                if (x_result(35 downto 33) /= "000") and (x_result(35 downto 33) /= "111") then
                    error <= not error;
                end if;
            end if;

            sum_result := sum_limit(x_reg, sum_b);
            if sum_to_lp='1' then
                lp_reg <= sum_result;
            end if;
            if sum_to_bp='1' then
                bp_reg <= sum_result;
            end if;
            
            sub_result := sub_limit(sub_a, sub_b);
            temp_reg   <= sub_result;
            if sub_to_hp='1' then
                hp_reg <= sub_result;
            end if;

            -- control part
            instruction <= (others => '0');
            if reset='1' then
                hp_reg <= (others => '0');            
                lp_reg <= (others => '0');            
                bp_reg <= (others => '0');            
                program_cnt <= 0;
            elsif program_cnt > c_program'length then
                if valid_in = '1' then
						  if cfg /= "000" or scale_cnt = 15 then 
							   scale_cnt <= 0;
                        program_cnt <= 0;
						  else
								scale_cnt <= scale_cnt + 1;
						  end if;
                end if;
            else
                program_cnt <= program_cnt + 1;
                if program_cnt < c_program'length then
                    instruction <= c_program(program_cnt);
                end if;
            end if;
            if program_cnt = c_program'length then
                valid_out <= '1';
            else
                valid_out <= '0';
            end if;
        end if;
    end process;

    high_pass <= hp_reg(21 downto 4);
    band_pass <= bp_reg(21 downto 4);
    low_pass  <= lp_reg(21 downto 4);
    error_out <= error;
end dsvf;
